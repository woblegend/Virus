MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���si��si��si�ld��si�Rich�si�                        PE  L ₆H        �   @  �      ,      P   @                     �    ��                               T� �      <�                                                                                                          .text         �     PEC2*O      `  �.rsrc    �      �   �                 ��6      pd�
A&��p�����B$%�����]^f���������&ؕf�X��Ж��⠕a�ݻ7L�������x�E���S�uA�qY�7����d�7�M$�"?�	h����؎��H���Q�н
�7h8Q���w�b�/	��%YF�]��dLe�7�d�XU2���"F�\X?3���`��;:�w'ꋎ�C�z�,����4@)_ǃfh��l�u����w��D�`� {#����-�,7��C"!�P�~u��}R�f�S��c��į@U�+^�Wڟ3-�s�n�3���(�����<��[�Yp���b\;�����:�(���T�d�}��<����x&k��	2d�d&���8U^�3���L�uв
�ٛ��1|�JA~�0�V�_�ɱi,�N�t�w���L�L�`$�M�
\�n��X;�S�������'9 ;���/�`d�3C����R�n�o)=2�XBk�u8pʏ�W]b��J#0��t�a�����Uۆ;�E�0�[�>{��Ru�JU%����C Pd�5    d�%    3��PECompact2 24A}��ᣜ�CN��NrS����x�-ܩ�/�%5\[�p�� �LC������k~N����̽���[)ݢ��8e���������3�����N�zs�Ր[�� ����������=�߱��D�h
��ZZ���g�h�XE����\��~�L�I����^��0#l�"�m���G|b�?肺�wT_%AN�~ ����������*��>���'��л���_�p��q�?����/'3���z���(3�UrUD�"��<�7�*3�T�[�����8����-�q�@�Z��L�J��&�ȵo��F�ѩ4j�T�UjlÑ�T�3[S ���ƭ�%@R��Gmj�H�b��E��$Y�_([h�A�v�X\#ցT���D���7:�����zǌ�3J�#T�j���Al�I���En�wZ#�|�oN6�%R9ȉ
`��@��Ҹo0a�' ��}��m�啗Y����R�{��J;��~����Zq��\��Y7Ǭ�D��n���"���5���E�`��kN��G��qyx�#gg�:�b.�H
D-�h�ĳpz�,1NQ�������M�k�&_���Ұ�Gk}���n���F ��4�I0�]S�4ߦ��nX�Ûz�da+
�:5�@��P�ʣ=��A����T�8��W�"��8_��"�]��s���l���iEbv�W�>�r�� � �}S��W%��(��a )�E�,�e�@nj��I��-$;�B��n����UPƸ����[�������ϖ��K_xv�ZV`����U����ؗ���$��?�P�p��o˻4�':-P1��αv��'�3*%��8���,
��J�.��4���F����� ��������&F�K�PdS��8�A��_�r��h��5RZo�
f1�	�-0��<eh����p1�>�3r�ǕA˕�w>��Z>��~�9��?{�#�*'@����ȕ�>d�Ѻ��>��7�-UW�#��ymI ȧùD�4�ŵ�aT�$�"��2 �$�ā��d������c�����r��?�p�	� މ�;J��[Ŷrm�D�-y��٫RM�@g,���lT��P+�Y�N~gQź��5�W����?�Y��A[`�SB]�Լ�xn�C�HI0�V�Y�f�l`����k4�Ee8�i�pF�BxE�퇘E}���e�f�̘��D�kCK�Q0T�'k���>ͱ8�ՍP�]ȴ�A�5�� ���i��o���bE#����^P�k�&ME���^D]^�c�66��&t���Q���iѷ9ȗ��g�Z�!�2���qF���l��R�К֟۵�� 2<UJ��u-�E��E�:a���~_�5AP��>V�lz鹭>����݉�?�A���E;��RR<ɰ0
��{n�!^|?�TY�� w� p_&�~�w�Z�%��EN�Os_�}u�IȀU�����U��fw(m[g�����M��9i/�%���:��O�q�L���
�f�7���ةl�߼@������G1�r-�_]���Q3��UhC~'=����"1b�/�gS@���I�D�����:û�}A������	u�oӱ��Z�G�ģ��#��zב��^���:ŨK�դ?7��؊�O`w������5�Q�R�9��af�ɣωs��ϊ�o�,�`��<���O�ǅ��s�#�BKޔs����� D�3�P�ek}��k���ɾ�+T8��'m�a(����r9�gl�d�X-G�aV*d�0�K_�����0��?�E���9;�UN��@V�Nz�iA����fY��c�������� �.]�8�� BK]!���`e�u8���	��� $F>6�-�����c�i֯�XK1��r�� l�n�pχ��|����d����J/��pc$���a��;�lnYr�f2+��c�yg ߙ�˟rǁG����w���`g�yy�::��[7V
`W{W�5iڃ�rHV�;��C�J����b���z,��%�
7s?��l��E�[hK]�"qT��wڊ��&����~�7��p����![��ĩ*�;��2<�c�L�*/�m�����~i7ǁY(���B9��*��{�Ģ�V����`N�3/�[��P{��h�b�zv��Π�<P��D�����9cD].�1���i���,��m?�ׁ0�=��к�ˀF������/�+KB1a5����ܱ������렪�n5[=϶�< t�����7)djlP��������HR�A�4/ <��j�F�?�S�5��W�ۺ
-4mI�؎L�6�`c�[�%z�������a����}�f��-F-�ӇU^w���ڽ���S1��~�)bB�,<1jK>�D������$�ҿ�a�c����	�bϰ�
�fV^��3�r1����ofvr���&)<�'���j�?�g��t�	R����}r �*�3���2��-/B{����d�q8]�De�1�#(Y�Ŗ�9ŕ����=�Y���O^T�Ծ9���_Fb`܏e��i�K��Q]�b�=�PE��;L���2>�G�35j�OT{��K���F]!�(�<���DsҐ�<;����J$�|����]�.1j�o�,�ez���;{������hv����Tm���:bKh���Q���ݷ�ډ]���9*�M��.I��D{�)pn��������Q�ih���5�y5���N>~'���be�����E�|}E`x|'�/o�k��v4�K?i����0qVS��$b�|��[�x#�O��v�w
�b�VQ�������[��v����昳�oP�7�ېfGA�\�t"�(
e'씝�� 9��0ܺ�������t|�W����2M��= v������m�4Xr���\Yy>rQ��qR"3@s����b�H�?�v�r�o\�5�y�V����Y��~e��G)8p���W��mG�)sO�N�%$8��o�߾���_I|����	*0��|�x�Q�]������c��4���93G�Gq���L���3����
���U���`��`�z�=���?7���]pж��eXG��]�R��0��pN��A�^mԅ����^��x(��A��!_��6�����6�C �N��F"7.q|?,u7"�sp�J�x:��ܥ���z��e�P5+��t�����󏾸fcċl���K��yK�v�!i��v!�K�MG�5Q��Da
J�l�C���"kq�܈h����"
%|[5�&o���4��������Ky ���+
��G�SY�뾢��?�ps�T��%��n��'"j����]{:�J��D $Wóq0�!Y�Jc/�I�'�R�n����j��P��A��X�	�[�s!
S�޷�Y����Q���dn>�Ǽ�t������di/���q��Q�>#5���B<��B�̼Vl��q��`=3 �f��`�eP��m��W<U/רŅ/�`�l
��/��ļ�'M :+/?�{؍���E����{y�*	)J63P���<��Zx�\V*���э\b7�����w��zb�*�ڡ���np�����'\�dU���KJ�́�K�G�o���N�"#��);�
��`s���Lҷ�Cd��o�J�9mOϵ��Ud�<��vU�/aJ�����*���v�C*�I(��H�{�##�������$�N���s;�ᙅ���q��w�ǘ��cL�qʜ��1�;��1ي�Ϋk�Nc�l;�O�%�*4C룸6�]��bM�j�uc/.�~�"A-g������$�\c�d�0u�u�u��|�5��n=�%�-X�j�s�g_>+L%�n>kLA,eēl����r*n��ǹ��+K��M:>���	�xSjF�Dd��"d�Z�Q�ju"��n�ϓ���H3�ع4������ ��B�:@/��hq�Cv$<�<�R��h�3�e�N��[�����+ϿB��\�-�z'5�|����|o+�a�Č��S[�@y��Z��Er]�+tg�!o��~r/�^�e����ҁ2@:a�����ִc�L�ĺg�;A|�F*�PW�Y�D�}]Q)0*�A��P&�R������@_��݄�>���?}eu����Ç��D���x&� ^b���0�U�`E���u^�-�
�y��4*���
du�
d=�17[KC���l~^qbz�.׮F٭cB��]��L]�?V��F$�լ�2,z��7�B�nĶN��B4���,Kc�; �}p�X��u�Gl�'<��<���b;����B���0�l�:�D�*e�����>�H碐��j��'	k΂H�]z;����x��6���dG��M9��UL���_����*�������.���o7c�]٬�1f$f%T������~��2<��b�~��Yb�t�{ccb�ԟAĥz�04x��K63�����<�����2[s���U�o�i�u�+�>A@u=�p}�󛫀e״���Z�f]�޺*c�����i0������-�=s�d��c�z2���_�+�7@�'��~p��s2�#��lpvz���h[����;$�cG�c���j^����I��������u�~zR�p��N�������.��ۡBq���Ź��D��Wb��.���R� �AK��аW�y�����؟B���Ⱦ�l�=������VY�Q�U!ƀ��7��@FBu�m�e��6ُ�D=ͲLQ�@�K�T� s��922�i���p����UtW��H������e�s
<d�=� {ڷ�4A���`��#�n/�q�����f�ۼm�Xԧ4�IQ����c��Jn�ؘ0eXy	�%���w�@�5�"R�7{HF� /��%��{r��_D!^5~�c��WV�K��-5[1����?*�T���8%�=�)9il;�H�U��j��`��7�A��IH>.^F^�.3���^!���u#x�M�V���^)�݅S����XczK�}�6k"L��F�|�#��J�e�!尥����o���N�t�)rrbW2RM~��8��d����MN*���<k���D�惶��8Aȋ�y<��`v��^`4b�I0+*Ë�~8�荫�I=�'Y��zy�`���uW�d!?��Cז��`M���<��0�'�&��˨QVR�����]�5y?��]�)TT�M;�6(�{!34w�4�����&�<�JB�hk�y��.+��,����3�#�>��{��F0�b�Z���,�p�8h=/�H.��@�F��8K�=�A���cYvw|�~���)sY��R��U��%����Be�'�3�_̐ÅGK�9ia�]��V�Y� V� X_��4i�]��Zg9`5-�d��elG�S¾�x,W9q�i�ɘ���a�oU5�ங�Q���,�\��ͦO~���?56��U������<���� K��z�zS�{��	���/5��>m��I�yf���U/y7	LQ$�^JѦA$�
y�n��I�"V0��|���ct����R�����-��z�K�{Z����j����0~^O�U0�y�,�T�ϼ��d\�sٝ�S�X��z��9���'�^k��TweL��7L��vI?���m���["���������[A>�s���/�b�x�R#�}�&{�;���58�6���� ���#���w�iiD��wR��V�M��� Z�+v	"�r����wf�e}�ϼN��=���j"���3���Y�k9caD�/.�
hmFD6��0���[EG*�B��膝��j�����\�½��4�74��=k��a�醚�):{�Ю��"���u�2�9�{�B�Ӈ^it쿳qG�R`���kvE>k�F�p���Ao:�c"���(���.9�/^���!��FY\,��K[������S�Yg<x��#2!�й�D�YZ���kDvM�H�'��\Lك~c��<�/m*ׄF��4��O7n�-�͵G,ޭ[������Ъ,�����t̖���6 Ѭ����@���S��M�ܽ�{6"xrg���6:V67��k���=�}��R��t�+�*T+�k��v�Fձ���y��Z��c=[�G�@��⠃v�4��Ֆ&~eT����X�#�t ���]Jg��+ԧ���VS~�(�;Y�@u�������1�U�����_(��4��l� ��.}�ML�f�� ��B��5xqc�O< E��Ph�Ě�[��H���-������C3n��*d'� �e��BrAB�|���Z'�oʭ�����#Y�����m�����JC_O��ͪ����q|p-�{��ɔ� V���.�6��6C����2��3{(�Bp@��Q;�
�^LZ�`��N���~aB�����v��酏/� ��c��b���u_n|W�c���U�ܵ�4c�^t�H�z��ن��?��e� 7�<��$YІ��9юd�4u��O�bn�+���)�-}ށ��#Ly*��:���t�X��O��9v��s��u�j�$.����L�5+�:ϐ3	&�3o+kY�p"Vm���uh�=��`G��Z}����`�ۺ i0�-�u���)8�������1N��ޜ��U���n�4��Z�]Ɨ(�YC!"�Bō.�ŕ*BX	E�b.�X`��{lI0V�Yz���6l=����y�X�����Ji Ċt�ۈ��i1��Q����ۙp� Re�řa��QHs ߕGP��S��5��M���.�XǕlv�]��^��I�,���{s�U��Tz��}��%M��{j����2�!9�5�Z��f(E��OzDQ5<��>�iuS#�q���w=�B�]j"�:���n��n���+!�E��?��N4�^iH���^��`������2w;�z��Ы�'Ȧ#�: �}��E��5��QI1�EE��e}��as9kd��\���	S��8�?���@;G�ޚ�C����	T-z-��8(΂`?E[EHu�U�A� �#f�V�fc��F5�(�k�S^�?5^zObn�K0�A�Mzᦕ2�]|�b��k��4�of�J��<�N�,���?0��P]&S,��yC�.WO\v��lK�,f	H	��]\���!�4�9{ͥÜ��U(���e+ZhEu�Wy�qK5R�$�����>���|��a0E�6���hߦ�����h����&7��
��q��1ܐ�&x�u�����'f�H(
*�����,
�¹[����{헳9�R���"���H�H���`��q9]:7��N\��Q+Q��;����{���� k��N�i�\t V��9�e���/e��>ɐ-���.p�L��=�g��r0�E�]#~�)�]A�S�J�;�6�d�\�`���i���8�vFG����X�߾NM{,�k�1�)�n�'�b���|p8�8�Rk�ƍF�+� �6���^��k���ps����ZUh��WzQ*h�)�Vr"�{��Bh^��/L-�Y��6�5�I�B.#A�$� �~a�" Ppb�s�lv7,�$8/��"�l������[� W�>����'���F�p^��~=~)txٵ �{�C��1�v'[��4� �./�l�AiD�r����hS��A�ے�T3�! �޶A��}���܅��t����HqGٯu:�`h���H��AM:�l 1�b��1����о|���#C�� �!���-v�ί��ګ��Q�f1bZ;�%
��l���`��\��60�dڬ�@:Κ�3��R��&���Сz�-C(ƪ)c�:D�f�}�Y�"؝lR��08�� S��Ei3?����I�A{�o?�O/=v��®�	^��Kt�o��WY�W0w>6k����P[\���]�jѱt�*�d��{���)�{�;��fW^t�SdG�կF�<��[��Gn����
ǓNoV�ʺ߭���`=��Z�G���8��&�l���|נը��Ú�$�8�EՌ����\ ��aA���%U��=�jc��-�T��1��߼E*�J����H�����V�]�"���&v�Emn�Ya"�L{�ț�݂0ϮaM�M��n
]���?�q�/��ƉP-�9������#�xe%F�V�bG3�foE��=Y��b������rA����w����JWoٿ���FkY�g�&%C���ٞ�u�D~�D�?=�$���GbU�y���q�a���:�?�`9�6�i�"OA�t�~H�:ӹؽ��n9��	|_���5<�[6�
��}H �)T�M&<�����"J�i��&�]�aF�����H�t���=����)�%�~���/G�L�e�;i����u1�sh�G��g�Vث�7ò��d��8�v�<����h�����_�dl�Ĉ��a�kg�F��iW�lX�8����AJ�w?��,&�a1f #O��9�x���N�3�(k�OmB�j�X1d>� �(��I	/fLX$���%�P<oGm��3��0�7?���(n�AOt�8�}.� =5��hV����I�d��z���(�\ɺ��5�v�ͮ	���RI��w�름����׎�`Sb�N`���A�d6���}х\;�n��oĆ���R��?�����2m�&��u2l��o�O�F�
�x;��Q@���!�U����ٟAk�T�|�9=�뵡�
c�W�#�$�߻�Z��f�o��E��!�P�f���/瑿X|g�"=�)�s��6��3z]n2����"���p~X-$�1)R �|��qg����)]�D��LO�G��ʑ6S�P�p�����C7��-/s�J�j���?m?;�xz�B�|���2��l����'˺o�l�>�f��ĳ>{�-ӲkQ�vt^e�������ե#���T�-�@w�$�@q͈T�נ�ك�����_'���kS�<`$fV�g-Ӝ��pۈ�:<�����O���	�� ���0Y��0f�J��!@
,�� �xfxÎ"�e��%��lE�[uҹ�T��ԏ��ɠyA���6Q�&[�U BA���T=���7<�1��^)_9�ڏ��{*���`t"@�#��B_�Y��E���J�����˭�OGx�V[~�2�����<�C����c-���f;c51:��y
$��n���G�1x�E���Q8U�8	�5�_ Z$xy(�����1Y��,Ů��?��}_;�HC��#�_N�@�T�W�D����a>�c�߫��aW>��}�Z �aIzF����3��7=��'���!<��L�T��X��[�bY�__���q2��ai��D�9�Ǘ���h�l�ȁ%�6vB {Hn؝��ٌ��,�8V�M�����zj�1$^�I���Ʊ^W-�PPG�;��a��9�(,��{g~�s�l���>
�ɭo]�s���Cy3l<�vI��T��f�rz�+@9vTl�~ 9��	^�g���^a��4=����?�bg�*re2��޲^y�ZGA�9Q�r�<z��="���k��p�(��"&���c�9�/�`���\����Ǽ>w*����g!��&&
)�me�1���(�xb��X���l��'�8~�V'w�LQ ���~2
�y<geBF��x+6c- )�σJ��|��������L��I�<{R�d
[��!��R��Z�n-�\�+��_26[!4aAū���)�M4�Q���0��P�"b�x[4��
e��C(��3�I\fk�� �DR;I�)͒b*��� Uߕ0���m}�r��̍�J�v��DX�<��Y@=���ZH���<���1��N��m�K)�g�t��E�"~�u8�{!��PQ(![|\O1�ET}ʊ0�x-��}�kܲ]��B0W��k�B(��FeWT��>
i~	�y<X2�4��!ܖ͓\年�' "/þ��f��_l��><B*�@��@�]3���<�,�2�[�����d�8B��X5�ʿ<A��/��<u�#!�Ê�k����d��t���B�V��Ey;��U����G�P�Ǡ@z�ͼ]�:h(�*�OBt��t�Z�Cj_���i.p�ė>I�`��[qc��v�|gҎ�h����?�C,��O�(ڣy����T���/u.���rԝhuZ�%ST=Al���5��\�̢dQ<�?�5��.��k0�HMn�'r�����ǖ�(ʸ�]d}�0^��u��~v�A�[D<P8��(YL<�e�Ьp���x-�@�/?=� �3�x�6e9D�za)0]�e"?��F	y/vD�a>8�8S܉u ��}��ߧ�8��!��Z�{����"�I\������a� =��yip��;d�!S�Y��<�JӬ��B'�zQA铮� S�
��_�㙸nP���C:�4	�:��ӪL�7y9&x:\#����Rk�l�'ٛ��+p;�wgO��+��f����]�
7�YXH�vs���#q"و��/s��X ӵ�/��8�	/Z����9;�|���`R4�cqj�6_]h����#g_Jbx俋�·�mӽ�
Qr�A5v�4�(��φ� j��LA���o�T�7���
se��Ⱙ#	����W��k�0ww�ʭ��ܝ�8b�ߟO���Y�+xW�=��ļ�4/@���@_O@E�o^d\�n^������7{��F�)��r�.�ҍ'���G�H�$!蓯g$�V���cd?V ���r�$>��z�l>I����W�k�z�g���v2��1Vo�'`b��d���2����Hu6������=�g��a|��*4�Q�r��J���bV|ŵ`�b�ɶ(����x��A�^p�C'�����^̑�$�Z�2\w5!.\����v�H>FЏ�#�bV��y�㜀`�n0�fXIC������Z��5E�c�
3C�lkBb�=��N;T�Y��N�z�>N����$z��^Ȼs韏#"ٻ;�4qG�o���9/��EwM�a�^Z���<�D���\f�a-�U��#΋�1�&G�#U��~EH����ϴ_�ը
K�]�*=+�`J:�}�Q�v�1����Ɔ�Hr�D��Tڴn~-��&�(�/����6�KL���Uw�po��(���/լC�<7#����?�X��/���G%�d����O7ް���UKo���!�~�ز����4�Z���m�K�`���	��,%��sC>�eE7.!��Z*~(��Kc#=�����"�)��AK> Ku u|b'8<b]��d���z�|��:�sފ]��DH	��F�7�@�$��Tty��Z�D檻l"j�wVy�*b���FM�������:��}+q�	�%CyRڇ�;9�a;H�Cĸ?����*I��Ϸſ�]��������Տp|�jU--}S����{�������^~�w��/]��zm�=��9�߭��2�&QF:a\���b���kLҼa�H @���D�׌nW�g�#xuI�)��,���U*����r*i�|������+bOZ���n`~�aa�����V�r$�ٚ�Z�t�9?)>k#���x"�}�D,Z�1�^E4ޅ�e��X,�Qn�t�fM�'Z�Z�54d�I��;`ti�ss��Ը���1�MB��=g�A{*�TN���Rd질�����>O�i��g��T|��D�fl�l��7�ܵ�g�F��]�d��l�u���?�GF��,?(z+9	�����g��V���X���g��|�}�C�2	�h��<8�x�Cp�~��S�Ȁ�s�Xf���hC�|����o���qP��%��x����N�9������uȽ:�W,jԯi��l�"������yo��'T������w*쉒������̶꒘j-�}.Y�<��A��ՙ�\�'���"]ҹuT�e�5����45�8�«�b�gi��uL9�nM���k�p��5n��N�ג�pb��6�^/����x^����}��M��ΛP#��m��֠#N�*A`���V��m�jҷ����@��~��]��O>�L���V��qu�	�/�����4�jPԀ	[�������T�3�F�k{��� =����W�ˉ$�a�Q�ͷ�k�w�Q�zT���*9���$8��{��y�c��D|��F�c���7��_�V!��SN���	>�:�W}r�N�פ�n�RVG=���8:��]��@=0P�:4����<D�)I��f61�£�������䑲r��)@^̷�=-IEp|��젻;h�w�c�i�%�7��.W4֘�v����Hȅ�\�V����:����GD���7Ow�M�`p��r$gYA���=:��}�	���9VH�����"Zad�%9Ah?� B`9�!�+��X�&�R�b����F9��|y�r��mA�*4�S�6B���0ৎ��Y�T�d)�h�)�V|���\�㇭M"��G��DW�s�萫�G�"�y�F��r��a���� �������ۜι?.�ԡY�������t���g\-BSU��O�Q���z��cYE@/E: z���o�����/��^��� <_���D������B5��YҞ��NW�;�`���X����O��F��N�zu{Bg���p�8t'��YR�w�F�mO����(������Aq������=8�Hb���������8�0�Ny�]_7�.�����I�������b��L���c��ӂݧSe\�ئ(��mb�L�4�G$B#rX��#�O�dZڛRA�t�՟ ����J��"XoO� ��ٍ�iԞ��철�:���,���V�c
��A�ja��m�H}�=a�~�r%�y�]���b���HK/��	� b�9��^�TQ*�����Y)p�����n��p
i��)�<���Cg���Ã��!�pwY���㍵�ŧ�f.Ѣp��|�e�M�B���p�!$�����IK�)�i��04%R��hk	�������'TbH,�����O�8���|�Y�LS��FY����d���.��@ �n �
�>�{"C�d^js"�7*B _�O�OI,�����m���+^��+'��}�Wچ7�L4�^�aƣ�`���If�"c��7�O-))�F;Pw�B�z���Ѐ�Z����3���[@��p�+��^8�����
���O�^0�-�_�� ,a�n⅔�b4�鯡'5�o�=�^Ot����t�u7�e��I'$�Yi�9�XgMo�/�������:�̧����bo ���`��E<��cٗ�R���d�1e.��J@�� V蒪
��	�_�Y`�\8��[Eq=�Vαy�OSBe�cR�b��b/Hx/1��>���ދ��1 �(��a�� x"Y�HU��ө0Lb0�՘n�]+���S�]����^X�z�\�cc�*1�;ɋwh�Q�)����e�S���'�݃��T��[���ZJ��&l�b�9'>���������B��.���M��?�C��h!�=��.~���k�j��Ω�L=jU����,q�ߜKjb^@w;nf����p�������(���`����ҭ5��m�����y��ҟ״Na�@p|Ga�.uIvbK�\��7iZvقy�2,��d�N�L
���E�|��l�8J�Ͳ��[����@�%�7��[��밳�N:�N�)!C�°O�Q�OR�	S��k�}��߱.�̀����O��"Bx�e䮲Z6G��S"�@����_i}2#��N���:˖��&���{L&v�s�!�q��ˇ����T-}N�W�q8���ɸnI����6�.oe��2��a��<=y��I�NEYąs��XY��U������A��*����Anq�.�R>5J�u����2���s�7�k}���G�׮x���� >ڕ�[ԊErĄ.��_���|�q,��6܊���~��W�1hs��f��_�3��@�����yɸ��"4��q��x����r܀k����s_���H-|č��
 �6�.~ȝ��~_rZ�ԕX�:Mh��$ �Ý(K̒�N&�('ƺ�F�7U���h��}/���u�h��kp��=�z2�%�f�Y.��fؓL ��.=Okq�l�M��ȕ�4	)�s���cl���Z@�M(��n���ڳ�(5�P�O�e�TuC���3������������G�~��p�!tحx$_�_�rQ����H�{(TK��Ü���&�/;��Z���޹�c�O7�5u1����7��W<Aֵ���6�䭡]�G!h(����'^�?��6
*��x�2�(����8(&p�=QQ�l����@��S%T����1i]�c<�v$�?	�(x~��w2ܛ�N�-DqTl�.��"܉�ݬ��g9���0��.X�t��=jj�b%�8Ɍìk��O|JuBNK�g���6����=��#��amq���R�A�x8_I@������^���H-D���>	J�v|>x�W>��Q��F��\��ʁo[kLĿ&N
C�bz�t�V��îy��^刟����N���>a��H�! �u�c�׵�y3�E��mM	j��X�7_a�t�f�d���F�D�1`RkY#����Q�%���Y�訠j��)s&"(�Ǳ���tM�D�_��wF�E�Q(yQ)�|��;>��dx{�O�G�@��H7�h�� �Ն�־3j�_�Jz�%���<}�@�.Ab1�Ÿ�L�F�W�Y�O����G�3�����9в�hh �_���Bx3�R�Ps�bsf��o�eӉ�6e3A�p1Cȁ�P���5b0�e"ٕ�
��A+޾�,Xr�])<�
���Hp<��a�{?��-��W�v�WBuL��g�r���k�6&��8*��'�?��[��4?,x�ҧ�bL��BG�)&��� ���E�&��?���	��t�����s��?y���y��AU?(��A�� P��o�+e��Ba������<p�S�B�΋�5<kU��s�$�8z3�v.X�;XB���׹����� �q�������@	Jm��|-��pׇ���lt-��=ir#!�����O�;x'��JN��.'���Y`��oν!^��F)XV�L�u�����a�3O����<�n��O]N)�TSҎ=C9��y諢�RV�Z��F^�,(�R��(�� �r��k�"�o(C���@����n[��TEH�+h����ś4�,}����d�۔���H��Z�o��n��H�0�����G��mQvS��Y\�'nd�%7��^�pYFM���ײ�x�-�*��(�뚰����f>|<"Kۨ;�}�ZtO�	#9��0���O�1|���i��(����,�J�l���g���m�G82�9ѣ��~�K�����<|�� �����>׵\&6���aO��N#<ę�UͤuE;	#���omm^ o���K�Աܢ]m������I>�\�¾����~-+���豘��}���uTH ��f/h���|�����am?�ۭ.X��✌<�ul�����>D��Bd:g��ymO ����w���)Fm�뭣%`w���\B�]�
���*�NZQm��=�cI���Zn~ի��`7�
0��Ǐhp2S�b �T���ڴ� 7��
�d'p#���k4iM��mB.'�����Վj�>|
h����T��Gd���}��DlD�01*f�e�\wy\" �����?Fp=8M�yg|�q�c7kϔoT�j	#7o=�F�'���HRtk%���a@SqV��D����:������ȉ��q��_Ő����LX�N�M�OW39/�Er�،�KI[��.ޮZI����Vo!٪�Vh����U�8b�ݸN�L���g��E|W+��FIJ� �\�u��\�e� ��R����q����H~��GYo��n��܎�ƫ�8ڍH�f�����or��X�R��@��ʂ��V��$ϭP>.:��?Vޏ�LU%4ί�`��6,����BT*��ղ��u�x�u'��p�a��<԰�E|F�H��G?�&�������}g`iQ?��Bm{�9˗�r��. �@�,)��2�.����Gݱ��j�;��ܷ���FO���Sb����y�6ӝ��ϓ�m~��Q,���m��-���aؐ}kF����5���	��z�|Ć��yRUS��� G 5);`t}���uS��4��Ǫ�p��9�}���Z5��K�H\B�u���JG��ܵ���XH�r&��Ŗ^���w� 7<�Y\�c5��!��	Yε�9n
9��NR�����.$�?j�x9��"BB{������v��}%H�d�!�X��C�N�Jvc��
��E5�T�Lֳ�z������A���J�&9^s�%��#A-�ڑ�q1}-���#kё�'WY���]<Ѓ��jL_�K�sp�2��-�W�+��-��j�7�	�����zd��f��n�tΟҹ�Im�=���4��|�{�mj�\�Վ�� �/3D������K&<��@K��#Add�k��.�%L�-C0Q��i��=���dP}��Z��.�:��&�"U� (�ǜg�aQ-rJ�SH����e�����U�a�R�Ϳ�ar�_H����*��ڏ�_��'V�LyF�T}����<F�ŷ=Y�ar\���Z8�B��d���H1�A�p3_����Z�P\�BT�Ҿ��$��`���r�k��+wǏ�լᡯ�>����+؀"
e-ӕX�����s5�����
{<4�b� �ty�WV�#��!�|�^�K���#R��B�|U�(t-��x-��wqG��d̗�4�x4
좦��}���6W���@M�bL`V&�
D�F���0�q<���Y�͚��=i����V4%u�+Dg)I;��*�3�@#O���N`�X�Y5�Q�$=���%���T$u��	�k�k�9;���������� �F�ѱO�Ze��6�C98���=υ��e��_�DRZ�FJ�g���c�!9����Adh%ѝ��7��ɗࡤ��{_�J�7!���g�,k���_)�I�B���32�I:��������ry*�z��ፊy=/����Y=�Y^�h�*���lO������|1���0ayU�%T��Ri�����m� �^��NB!���f���X�L��4$A_��A��T`�BZ�O�4�Y,n*֏�`��KŘF\p)>HP�v������.�Fy����,U�t��**w(FG #�ꎄT	���z ��uTT��k��d��e1��(�6��bՈ���1wְG\'�*wB ����v ��+�x�
M���>�Վqn�9n�K)u"�r�&B/5#�軈���o��[d-۟ Ehː��
s��\	��0�~H��ռ	m��9^ӥs�2��ت��JO}�h>{���a����`�9՛S�ܬF�[�C��3�,����ӭb�hҬ�B���fY�(��^M>;���X[��f>����l��_����9f�������N�l�8�#��\�%�$�9�����9+zm�Y��W]-ө2��^)蕼��5�.(4��Cy?GO���ع�����I��.��A�ѕ�%i��m�?���".��g��S�����c[�#���z�7*:��]LM{
7Pˍ��;��"B`��=o*����O�U�	���x�X�Ga2b���6K�ZˑH���^`ڗ����f^[�bF�ϝ�El]�$���$����r��5R�XE��nߗH��D���.0UV�31����2PM���q�Z1�ܠ|�83U�f�ȡ~ ��7aHi�<#<�;��~��e�6� k���8+��X|�VX:t��P��Txg!����i��J��[��@�M* �'�>�::j8�0�61N���t��6�+�#�S>ʡM,��U�oq3�j�KB�C~fV��n�e��q��
��dec�§����M���L xF��e�di��7%h%���H��s?^Y�8`+���32ⶃ���i�?Ho�a���!�e1�H��ک�Aw��f dqx���B��~i=�C�B%�cVz�e������qT� w��k#�ح�܍�<��a��VD�	�3����)�B���[MC�}հg�������@�9����n:��=Q�x>d*��\�%?������3�؅��m�z���솴|�"��W0����F�i�mghIZ݄#�|�ԑ�,_8Y���Q|`��<^�2�[����T��`8r@\��r@�d�eCcײ5V�(�m����3w6\��J_�4(����Z�}��=�K(a���+��jpvD=-N��n���n)=�l��>q�\~zJb�O���ٛ|���vk8_&��||��O��?jըC�B��K?!%��nV/QDq�o����혀�n�E>kۢ��]���4���l���1	Yg��5v|W��D���Ȃ9ϛW>]������FQ��c�ٚ�F,Yk~k��;�����?�S'	��g�t/�׹��O��Qn�m�=��A�00O;x��x 
���h;S�^��mk;�)���
!��P�V%���>���OuJf"��)O�;ս�}�&���UKƈZ��Ƣ��
d ��A��󢰋&M������?�o���f�y���깛+����h�
��*p<�8׊\�(���2
ݣV>���n�$A��xU�J0���2�F[��s�b�������0��A��_�x$���G&�֎ ���
��=���i�#�t3���aW��Џn�5��.T��(�(�ՃU}���r�5z�콖|���I'-5W_
%���47݆kG��)�l��[��^}�%��l��jP��VOMoa�A�g��k�Ť�.�ld#�p��>�g��O��~	����W����t��C�����[l�=���$�lB�ň�!Zw��/��N����ȋ1� >�G�Q��$��w}-�B0�g��~<ܢ:2x�0P�����#�i?� MD��,�KvS�w��p�\�������k��9{�d}У�`�w}�[�9x�/��v�o,�m�	zjw��(m<l����J��z���$�s$$�'<a�!���(Ul��e9�xm �<����@��q�tn���CC讎�����K�'9^�.���l�L<(:�{cn�fOoU�հJ
���\a3�@�9z�� ���v��qY�]��Wm�&��F1�tH�6 W�6蝂'6G�ZpQgkV$Υ�~�� ?���!B��+�Sȉ#��l��3s���g͂���о���Ҍ��%�Oé�[�vKW��G��8���#BI��)?v2](o#�[mD%Y6pk����i;6���4��IJ�}8|fe���s�y���W�v�� ��(Մw�%e b<���c��AW��"�hU�e1��/��R�t��B��t�����6R�<�ul��a��1�U��i����m0G�4�k�o�f�y�q��3U�ݔ�ϗ%=�H����=U��w�XGe�EY=�l%q���P�����/����i��oF8��ؒv���/�Y����j�B���_A,���+f��p��Խ��q��Y��;�f��s4eW�����v��o)c���y����mř ���������O�Aj�BY�v�q��d@�G�E����� h��l���B��s��د�S��݃��������O�yx��)�P;�X�����"���|3�#�[4�]K��B͚��E��`7B;B��n��'Kjo��.����~���w��]"J�ۋ�cԆ�e��F�fu9U*h�G�p�2�|�k������z k�tD=9��AB�!1\1ߗ2�Q�(��s��uw7x�i�o��K-�~W�h�Iơ���n)R��gc����Q�}a����P�wF�GL�j�䑻�Z��-���-Ha��qq_�Ӳ�����T� X�qЭ��c�9���<�^�%b'���er������� �,���+gTX���c���5U+�P|h����x�ks̼Q�b�B����zۮDN��P����V:�B����:�bb��`���vF"�M"�>{UHAo[����'�u���w�g �	K�Y��2yBl���~U�G����)R���}��7�C[`"R�Ͻ�kw�ۄz�������܃y��w��KgG�d�������d�H���V�F-�K����M�+(}}��=��e@��O��?>W�rIad!`��4�2����r�\+��V\v'%�}c��{<� ɕ���m��/�c,pP�c���x��u��J@�x�fo)�TĠ�FfH-��胖�3�7�>�� w֤I�%g�[;����Y������ǔ�E[nY�c�r���K{Q=PG@�ޒ���v�<5�
k�ί��Iع&1��ļ�;T��9��A�	�P�ϣ��Q<�95�c�J��@��״c��t�mR���U��.MR�co}{^�L�-�;P�ɥ'�7n���E�(�P&bǩ��=[���橄<	�K�/�!�+���#�me�*�*�j
!�z��inf]
 �uT�n�D!���;ax��ڰ�#��fC���@0��;1��hή^Y����0��7{�}2
��
�d����\y�j���Z�kT��2c����r�QN����s��N�!��F��v�Ku�R�0�/9�$��a>/�ƻ-� ����'�AV.�ʄs�Cv-��7g5?{��"�	F�#G��
Q�y�0s��9�1v�&!$2�/J��u"��0mAQ�|���w�H/%]Ɋ�Ay��a7��֏h��m����_b>(V~\)9p\��7����(��Wq�E���1˳���M�T~0r7�q���=����:(kX����|]�i�5^��b� ����b!W�°O�}YS�*FY�2��ըDO��0�v0�d��K����,|{��m�b�;�$�����^�%�Ƹ��:��V:g�`g�����6�w��|JXO��g��-���ᛗu�к�)4ؽs*��N.T��SJ�z&�߳yUUuk��?�'��
S���Xi�N���~`|ҩӢ�
��z��nr��^u���Q��R�����VQ@�k�|��JX�&��5��Z�Z���O��;���P��@F]�AQp!Lv�����;��������a�Qr�'��1X�F.�1$�+@r�HRo�Rs&i�#�����j��NQZ�M��5�ь+��?�B!�F�עSƘ�O��Wd"t�j�g+P��+����I��fu�ay�3�_�p3���0F��Z�9;��d�'��j'�T�5h�Z���Y2i��*��|�U���'�Y���(ك+ޔ����2��x�V�t�) �HZ��-�L;�ƫ�Qw�[�oW.��*��GKK��^�SBj-1�H�Gt����";�%\V��N�|�]'����=W=��%:_��n�"w���_F����tn.�瞀�Ѯ�L�=�$��8�	)9��[Q/���ɗ+�p��8bj]���6�/�[۰�����	#�;��W��o(�>B��w����A:�"���̏Pϸ�.���T
H�ͨr�^#�{W�BP�
�=�[H��U�3�;?�j�Ik�D쾇B��[i�>���!�9��h��U����v���t���m�W�
D�}�3$f���P�>���"���u�'����3��6�i�� /�ay��*x2]�vZ�H��ʙe��$R�1E��Wi�$3(�Y�ṯ\�����ʼK�4֓g7)Jt�����QC�i���!��<��G�ߘA����Bs�e" vם��9�$;��;�{������x 琭���t�=�I�Nې������1��*��o ��^���5 �;B[f
E����ؿ��ݖ{��q���E_&��9�2�蜉O6��I�N�1ϐ�T8���u���i��>��xL�c��;��6u6�g�@��5j�4�>�-Tm)ܖ�1��P2����Bs���d�5�'��⋁ə�{al�Ե,���	�'�#�;��eM9���� ���h5t#��/�I�M$��/Rlh�C$�+*Gp!��~���f</3VC-�W$�)�A ����Vjb��D�3�H�{�3����D}s�9�^f�eG�p����v�����1����:qZN�Z.~ҙ^���"u.����A>V����Ȗ#��ڢDέ�-���I�T�Y�_*���9H38��$�>[��$t����b�����ODRd=���e��e"�l^�i���_��Rw�l�Ïc�b}��{��� �	��u!�1��{��F���/����D�<1 B�9^�b�V��S��Q�4�T��A� ��@1�~lA�6��������E�Wv�I� 4�ִ�MC�.Yp}[)��x��{�G</����O��)g�y�� �JKp��	]�u�X�e.�z9
����`v2�A�o.�����Ǥ��?�|�e2���������`�PW�H��$�9�p�G�@�x8�
�W�KLUo!?yK��/��󨷫����;���X��.&Ϩ��ra�����<)`�0|eS
�
đ����XY�OHw�����*Pc<X\.?�Bl޽޾gz�%{X��QN�Y;(K$Ŗa�9�g�����f�s9�S�+3�Z�]�}snH���[��l�s�OÇ�@G�9��1+�1EA�P�0a�$(&�˞���]YZ� b���TV��Vf�xE�|�jo5/�G&8�Y���S�G,R�A!���9���3g,Z�&ZZ$x����h*�Z�P�lwaա�MIR!,X����s��������GL:~��?��TDU*U�C��&0��G2��q��`の�y�P�B5��&�|�Е�0¼������ma��ܐ1�-��H#�����i�kZr&�2G�4`0-ΫM���@��G�xv��|��v�e!��JD�@1�����ȑ����˦���Tq��)���t���+�l��{�����7��8�( ]Ut�&33�*���ϼ��r�f�mU/�F8m����s�Z�ڝ'�D����slrE�jR�T6�XMa�7�\�7�\�LKA�6W�:��A@9���)e����A �r�^"$�x�׮GEz��XQ=-����,���h�6�D��lZ@������b�����Ì���0���u,��d&�d 2 b��d�U
�/���Yo:���o������u�
8_��칿l�:��;�q��";���m�N�� <����"��9����۬���8�nl���d��T�\�YF`bk�c��|ГQXe>�N��_|3�T���p����29M�����&�	'�
'��7z*n����:,o�/��H�æ}����3�ۙH�F��0�0�(Y�O��(z�6ț����Y���*��#C�Z���+-������or��I��2���Ns�lu������3�e3 �-6�����g���+�]�����-�!�2d6�,��}#0F P7+I{ &��pp��Ķƅ�Q��8�q��4\��S=l�����,��*��2�lK���R#� "�YD]�S4�<�j%���@M��Je�)s̀�8���D����:�C3��*��{z	�y�C����4�钎�D����J��Ð�Ǳ�4$�!Ͱ~CZ�uM�)< ���A���x����9�kju���ЁKؔatt��/�Cx4��|�}�.����$�U��x?�U��<�3{����"T���Qw���L�Su�=l�g�3���ݶ÷��^��� GE�B��| �J#�q>e���r9Y
��e�Yf��K������$=뫅�ppxx�	�����B�y��|}��!�8�r�v�]!M�>R�>\6�L\��r�vb�3��ݮ�t0[~��2�i��#��'{�I(4���􃱚/�� $�č'5�G���Q��8vMPOJ8HS>�=���=���}M���8:��U���O�,kql���v��I_Y�lX^�Z��y�$�_��IH���2R���W��)����q�)�*J��J%s]g�݊AG5��$L��r~�����Ɠ�H��C�%�<o����������v�Z����Lf>��퇙��cٌ-A�vR��s`�r��Ps��39XU��?'�*�>��ۅ����_�� 9�d�^N�Rr��,|�A����:�V1@���a�3��!I'�)��yGu�����5�(9
\&�M�ޯ�{�s�2��X�0 Ӯ�y�!r��d��>�y{7��?"��6W/?�z��(Z�ʁ�IL�Y^���s3&����0ʢ�u�.Z��t�E�&�ݙtƣ�,.��}oy�[�^a�1�;�YR���H�ey��[��l�pWnu=b[�1K��h��\*ja������<��i��eo��o���V̽9IE���<:#�.8�����ӖA��e?�CW�;:����H^7J��������G<��w�o}R�
�|��tr9�צ�\B}9T�;����E���P%q�� 1�Hhӕ*��狐]�@H�4yi��3���U��ͷnx/�c�Mm��gM�j�_�z�>� UD,�sK^a�aLU�n�+V�c�z�J�|��->d�`��kZ�A�v�YY��<%�b��r�p�d8����9�h/#��j�[��!)?$Oe��ڬ�c��O��5=����bp��=��D૑[uHY�b�R���:�L֗����˷v����yJ�ɸ�(�"�q�����-�|u��� '<(���3`�&N5$��$l�96Dfy�>��+U��&���FT� m,����Q��MӊiK(�x@��c��e��W6m�.��՝V�(����1��we�;���P]\���wϏ2���	��X�;bΕY��"'S�èX�x�-�ި+[��[ P�?�q�e5�:T�Zzޭi�������S1]܊}�%l<�|*ۀ�{�W����[1/3m{�`�")XÁ�%N��&�m.�О�g����`�`<��M�ǟ�K�w��Q� y:ƸYM��R�K&5�0ԩ����R/���Њs2�N���q�z�D������I@�S�,����A�S>�5����̵��,�
D�¹�K���:�S}&e�����e�_*@��nC������*��Nky��*da�FQ�Նz����[���n���T��V`�ˈ�}8�ec@�(u�dn�V�j�~ZoH�������v��X%�x$���Y�r]0�>R�E������ ����="�U<&=a(��f����=bY�>�:��$��dW��aw]�mDwFJ}�O�͙��j�Ӿ����3�|L�Vі=�ڊ"��V�{�u��4�z'qAJ�L���_��g��a��i�J�J?�`�`�/��e*��?��H�G��I�P�~��d�� X7�9bKk�(�කy��r�p	���ˤ���ma(i��M#�Xq&���|�qq`��)Pu�J�~H�e@r��ޡ�l��8'->�rf����%�n9�"�gf�J���<�wXfr��X.-���b�.������ ,��O��aMt$� l���"q�l��+�^=���;'����T��]�(�N��Κ'��(tX��c�����O<��_�+�I��8���<-u�Q��OQ�4��p}�ѵ5�f.�;T|���Ǣ��MB�����������`ds��P=R={>Z2!�ί�M~�݇i-%��>���� ��&�jwQi�4P�	���MOQƠ[�-�V݆�!�ĪY���ƕ�<���^H�'�I���_k��Qq*�=4As$3�`�4��i�wɑ�T�g�{M�3}�j߀$��G���yu�r�,Ԗ�T=U�ӵ�a�ot���&B�����$�\�������M^㪩i{:%�T��צ�Y��&�?��,SP(%M�+e�b�j�HB��DW���������=J��$zZ/���7��h�ߴ8���I�j�H.�w�A�k���_N}x����c����X��b�Q�=�d�-���iϚĉ�n��I��჏�\���+�����9��W{�KA���^�V��:-�Qĸ�^d�Ot��x)4K��@=��s��<��ܙ'&/V�U����$1	��e4��B�y�ϥ�b �m+�[Ѥ�'����נ�F�m��W���&/�z�z��W�aB׻�zǆ��L7�T���v�4���q �pp�+���sZt�"v�F'#:�����(Λ`\���k�F�oѪϕ\��fpXr.Ow���(�Dk�yI��|,�:�Qi��n-�~�-�r��b;��zl����/�A�|#�0����g�]�h��
��7�{W
\�7�x$� 3�:�Q�G�=`띥�*-,�k������A�`�:��f�j�(F��`^�!NNR,h��o��q��<��<8�ɣ\jןY&�h
g���b���^ʋ߬��B�=c�����c"L��l��$n$m�T���4_-4���i����f>aJ��<hwp��.9IR��j�̈́��I��K�<��'?�f��[��Cd���9���7�r͕�ک�A�?��0Ǫc��(��"}+�e��JX0�`1�N�j��
�����l�|Vg�l�G|�}|������°c� ;�O�-m�Ξ(��9(F���(I����Ӗ\n��<�ӂ����x2Z�m�9ؙ��L��dDA3	��B��dF�J�%O@����K�妲32��1Ӄ6�<D��,�HUL���XW!��ɷ��t1�ϱ&#�gp�� A����~n�9׿�7���l���?�c��`f��K�����,Rm.v��z6�amk~~��	q⬁ٿ�NA3E��%����h鞌kT�<�Ou�B!�eK��t*j�|�RN�`e�����{Ԟ=�ʈ,)�y�<1���������J�k���<����1���G��r��Q�U��oS�:���d�D|Nk��F��ݨYm<���*a�R#8�:騞[0��k�.��k�36�(�x^�j�3��bx79�pQ~܀�K���#�cz��ڤ].L�y�������\��]�:o�EaL#!{�c��0jz:|pV��*]z���Zr�y�m�=[>��K�c�>U�qZFn5�D~�m^������FU�V-�/v-���+�{T�qc�A�3O�WEhx����U;�F���`���V�j�ȓ�:?k��A��uC��|!���;&��$k���*v�	�w(���wk&6�`�:��3F���0��#V�u�A��[V����Α�v�G�����$ʩ���f#&�}N���#e������WNjMetļ���}2%��������ס'H{7�gۑ)/��C'����nhR�ahTUЏ��v䭐�@��J/��[:0��y�]K:���Z�w>x끱�g������[��Nd%W
&�4�<�;|�b�(,*���Wn�5�y��U�ᕉy�J(���������we��׫R;^D��s1DQa�>�4���������iEc5T�\��ͦ�*H��A�B�XVK���2�~^�'�+h�����>�� l,��#{��UfBvi���]AY���wd��Վi������)�Q�;��3�`�:� �,uHx�������#��iW����C{�}K�st?�ubG�0�{�,�R��'%#˯� QS�`Yq�� -S��!b�v�J1�ڶ��h��W�ޏ�	�v{P��?��e`��z^����)RI��o$<� {�5};�mJ�W�Y���� ݡri׷;I��x{�x-k4P9�����?�����У�|�3��v����՝�7�����u[݋�������}�D l��в}��P��R���"��.H��,Q�
�a6�4s�ZX���R�Ƨ�b�����t�ȣK����r|ͳf����L�8��¯��H���_d���;����f�Xt\`�q��9���sL��SOX��ێ>��/԰�,�t7+�����"(�޵�N�{��G6#K��Rr
r�Y���u�͞Ip^/z�^�15Z�Sf�5�}�]�\�!MTZHC�M/���Z0 ���}��T�f��&�����8Wo|�������6jP5\����cZ�H�����k/���y��掄�a��ތB�m��TD(�I� �����U2^����t���N�T-�X9��l��y�H����r��zXC�PxD��,��n�9xk�a���JE���|�3U�1��{
��{qɄ�eI��f
�nCL콳Yt$8�(u�V��jr���^1Cq)J����\8��=?jC=���!�ў�-=�\���.+��>+)�<ru:>�]�)��(�ƫ A�;�b/[	oҶ)�=]4^Y@7�C�}����'A��E��dt�;���\�B5�[��ՕG18P���?zW�j���]��،���I:�	��/	%@����r ����/��,?sz�O?����=���`ZU?��ұ��mO=g7z������1�D\�1�p���X�J�il��O��v��U�
�ד�H.W�ۚ�R|�s�x�Rl����Z�w��)���t;Rx�e��~��3ioO�/{�h>K����9Ï<�n#��T�;y���Z�=z_p�j����{����ѳ�A4F��y�7F��(�cщe`-�I�\�A��.�}W��RQUԏ.��ߩA��.x�����j�nq��`�I�_qx����f�DX�֥�����{�q
�~8�]�����;R-y�iG_�v� ������Ý�Jp0y�aB�ǔ��F������qhΒHO�v�E�<ȷ�n�'�v,/�"��G��o�������(���%Df��kdFFHBk߂\�fR�S��5(۹�X+������iO����M�?Ӹ�a)���=㞁��t�Q���M6�!����FW\pd'W5q�^�\��@)�r�20������7⹆�[bš ��+�1~�}e&z�� ��דL����E��])i��\�J���Qw&���ʛ	cF�v���=����Ɖ+z('DV�������\��<(F���(%]cE�ֿ�r�-�}Ȝ���N��=f�� �s�Ew��1�ow�j�{����ƨ|�[R��?�Ж�x'��#z{�cʽF�#�_i����#6�R��t ���D�rf���e�W�@���O�����<L?��N�`��d��w����$?$U&Gl�L\��2�~��'1���{
쟂=�L���gN�L<vE��`�I�5G;����_j5��_57�^5ؔ�CBP{a��|�r;������h���S�O��=�;�~��R�W����C����\2��:~Z]#  ��΅��\0�0'�g+��_,@�
�D�/�C�3Ņ� P������� Tw�=�K�����\���ϓhor|{��^�?��l|Wp�����~�9°�42�[�(�E�%�	�~�i�?�%�G�qSҎ���Çn��'�������c� �a�$�s�����$�M^$���R�
F�#]�1{ǋ��n9�~��Sۭ��[ÁC$�P����X�"�/����Bδ	�~˦Џ�&���,ʨq���$���4]{"�)��/�� ����C�mҚ�*~�1��r����� T�d�ſ�v��O��?A���y����\_��oӲy�"�՝c����X�LuL�T�%	U�ҏ�S�e�j�ʨ�v/^�&���m�dv��Mσ�b�9�?���h�����W��J_@����r4�=	�,��q6�}n�;��5�SJ{��/�TuMan���a6q��"�~�\���F�K�g�c�BGj�zu��V��K[E8�ør�i�/��V�*��\�@�3�r��o��M/�%W6�l�B������/;|������B*~���_	�K�QE�O0���ln����@ŗl;��ɇ�S���?K���)�7Q�'?����0z&�#��@��5Za�{�u��D���������>��7>�R�T�X#�(��L�f�*oN�Fm���Cu�
�Y���eq4�рO�O�v�Wrթ���ᆺP�|T�zu�d>8*�J�*�A?�9j=�wPG|�~���������'|]8Q�^�Q	iŷ}�{ آ�kO'n�_�|`���yxrr��/��a�&;9�C�a"n-.C�!x|��o?b��8�K,���\4�
��dN~���T�{�(ug�ɲk�%n��8����0V$R��{3�ф>4#�]F,�Ə2������6[�l��_�dm���oY.T�=��G�P�\��2�����,.�#0N/[����l>��N�!�.`�B��RJ3"b�X�hK�^�sd=ڭ��S����h�Tn㩉h"�D����n���+���:�-@�	x8�P�6��xO�%X	Y ��R����*�*��9�Y��G�-
���3`EpK�X��#�tbW��WB��&����:t��c��.-����8a�!RRQA�05!Hwf��l�̟e,M�	�v�+TP}˗��Nc�V��u]�������^{dOiN��E���çd��$��F�S��p����h�A���Đ��n�e"�Ru䙗�9�3���M�>�>��X�e��+��2o:�Fzm:-.�����v�'=��`U���9��ճ�gsE1:W�ifS|�]��j�?-����2N����2�"Jĩ��Hզ�����[�����=�{0kb�޹t�F� ��J�� ��u�LpD���/��]%�7W��R/v[՛L)���*Ze�#O���и�m���D��ه����M�q�S��F	���*�%�s�Rǎ�O}��$뇀�"aqb�'6���ޕ�=s�����@��v]2Z��g$rࣥg�����:��0��	����5o{�8��j�k�]b�V��g׌�'���.ѨDzKL+?�����Cw�P��a�:�*l"H�&sL� A�9�|c}���w����U�ˁk�N|Cd3b5G	i���;ʂH�`;�����z?32J�T�}9�̗��	�,��N!m���~��[��]I�c&k}nGe��>ĩ���X���u�C0�)��3֬����g����mX����a����@�?�K��A*����EpQG@S�Y��H������O�Wި��߆Y?�o:�db�z���U�)�l�_�򓼧�_枩�%��<4�vea��$��w/q�>ߔ��e_���x�ǉ���<w������I�P-ee���th�e�p����N�XE�(�3�Y9gL�Cw#)�����_�B�z 3D�Ϝjc%���r/T<?�>�"����dffI������e�m�5������1���=U�N���n�w.��2�y8�����Ǩ�P|qN��y��@��8Pͽ��E%A�=B,���T��ԺF���Ŝ�ޏ��5o�0ҤM��kf����M���uӴ��;A/�T#ٲ1���ka�敺@����}����=g~�.P�_s�΅;���`G��Υc�e��$��f��'4��Q�*����ٕ��z�T`��9�j,��Db6��C�K����8����\����H�Љ�07nW	�,s�|5"!���q"u����OT8�w�b���0J;X1��3��|5�~�����Df�y��?x@^f)�ɵ]�Cg���L��w&*X '���c��J�x,��s��,�Ui��S���c�ϜMOA�G^�y`5�s*��~-o0��)ޞ�z��ݼ�������}1�A^�-S���W�������kBV�����+�Aɦ�K�g4/u$+��<3�� ��i��8����m��aؖ���;����NRT� p���$,���?�}���,�;r�4}E��іFhcR�{�H_� m�b�s�&:(:�yt(kL�����4B�Ʀ�Z�#�!y�����'�j}���_6��wn�C�9I�_��t�0���\M%�nX?�@t�<{�lH�Y�q�

	���qWk��>�w3���B,[���ՁR�7����Uz�BI�Z�f;4��pBH)J�a�G*GΤ$�ό�9!�f��]w5�z���jN�6�|em�c�9|#&b�C���8��Jv3�z�`]vc.��N�Q��6I��g�Ƀ�d�ؓ��c�?�� D뉬��w%��[bH�7T��	.��(�����4��9L�e�ғꟃ����)b���q��
6��� ~1䦆���8��w��o.�gj[f�ݝ��
6������<��k��(��Ӂ�� �*CC��rJ��-��?�jU����J7����������7� 1n��p |{�F���QP�����Pi���d�Ԏ��^��k�i�7�&U᪕��|�7�k�^����[����l��� ����Ȣ J%[L�h{t�����Wbu�\,t��/"J�N�d��	���ی���
Q���)�f� g�����:yii��f,V����3b��[��'oZ��N.� e$lKV��?�p���P���S ������LB�-2�����nA��;h��XZ���<��S?�Fkd�'4
Vu%M�ɒ務[���C�,.�Í��լv�ǐ_p�+3��;�f��D����"�$��	FF� �ѝ��Fi;�%�F�2Ϧe%���!t�)�7�I���4]*�hU0�.K�-�hF,�;�*��+T0�e�%Ϭ�{���dտ�Ǖ�����Z�ed0f�&���~�^�����{��
*�s|Bi/[�q��],�Z��s}��=CO��7��g�?F_']9��2�2�0z-�^�(�=K�rˎ��F�c�br���7N	��Hɱh�߫u�����.�CQ��\�M� B���̱ɦ�|��Rq�����z�����kB�9�97/��̩���	�5J�[PJ����b����6��*�8jC|�r6�ox����/��6i���e���V����Օ���T��6��گ��s��t��P�M��E�-�<�,Y�U&�U\N�>�@�U[�5��\sqW�6�[u�����s%n;e{��o87&�e>���
��O�6�4c��!�eO����	�]��N_L��X�K�F�>d+ ���Ǚ�9E]��8΄އ2YH�JX\��#���7A;������\K�٠[�L?_ק����W���7��9��ZBZF'��H>R���R8�<@�_)A+U����ch��Z��tɁr`� =�f�(���f���[pR`{�A�i�N�08;�|uԑ6�yt�yR8�ho.�.���r9���.X����F��x@�:z&5<m�aY��8�\�;��b<��v�c��QֹdQm%h�� ���(Ee�4@7��#H�:"s���@"�y���Փ��f:-�K���Vl��f��������xf�gi�[��X;n?�A炯'l�2�\����@h���ORM"W1(#�	G� RFm�5朢�uF��I�x}���v�Ƀ%1
(�&��f��캅�%l"�� i���by{��Q�Ԧ��6��]iFI8�"�lA\H�N/�=���@"���.��H����~YD%YJa���ܦi:����w�r����*��+Rd���E��C�u��0�J.�ז�ߚ)1�$����±��
�j�g5ȟ�E"�?)7�}��t����1���hΎ6���	�(RaY�5�e=/�_��,w|�����r�x4(4�$C
_��~�W��W^�k.�C�.Uzyq��1Tpn��.���X\=T�O�0���jn�(�IW��Lk[]�d}X�MM�
��e����ՋT%�
�f��tl�����28��
��>���v$��S�G��L��D2j���}��w)�Պ�:�D����xqVIe����t�6�����dz�i�{��p���gh�)G7�\I�[X#5U6���yr=�-�bZ"~�`@n�8������/\�z�?~(6x�!��f�K*�'V6�P��sS&�*��<tZ	�4�E�\ʿH�zhpz%��U�%��푝V%�?���J��M݆
H�j\�¹�cDD�	�~ � ���|K^3�vj}�����q�u��c&��C��]�g�yO]'z��V6�@�%ż)�tuK�1\!��d6M�Ɇ�rI}���x�N U�t���7��7��_��+�F!ؔ���Io��fr;�ُ��b �E�U�F�����5I�h��mG�D0���V�g��ţR�3,!�GJ�|0��Hf̼$8��7n�;k�/'�c�}���=��a�H��k,�v���P_�a�|��{|��;��|�����B�P2�bD���Ğf�YP���|?���9�x��mP���>�N=��@�~r;��ΐȫ���Tb�$.��t�ǿ4&��`���q��\i�P�xC��I��-r�� ��6�?��1��9`�#c������?��׫���@ȱ�^�!�k��گ�'�Y����7�nҒz|2d�D^�M��\H1s���~�^���$b�� �V�)����s셅�Ë�'����:y��hCf�F���a@u��F׽\h\�q,b��*�*k�	��l�W�a0}E�m��f~�ǖ�6�m3u,���1�� ,��[��x��~�P�F�
*��+Y!��$�d���b�:��'J���<k���5P��O��L�ju�=WP.�a�#�GW}�_i����1k;�(XM�����}�ϋ���Sғ��?q�qh��
�g;DJ�o]Z���Ԅ�@,�R��F�w^Q'�����ZP ��ƨ��Y�wM�w����4��'�q��L��u:���Ũק��7`�j��X�k��y�&�mI�=� �~����*HzK���;|#�����.��tf��KnX���ǥ�K���KT�����y����Q�.Fs�椏��]�:u�Y���E��P�L���� ��hQ�����5�1Ç6��T�}���o!�m�5��H@-�gj����V�z#5L&��,�y�(���c���i�#��,Hr6&�x�>�������(z���S����Ut;�����ZkM�Gn�ů��%����{��(�#��G��1�Y������#�-��E��FID�V����A+?��'N��6�g&�3x�f�!��hU\�!Ӳ��ys�	�9��9M��n�y��je������[���g#�����qV%М�GA����!֭xҐN��j��ڍ�i�1��w�e,-�Vq�"�-���a&d�U&���t��OE$���Ÿ;!LyC�+i(�}�v�@H\�;�Ͻ��R�X]K&$�w�*
?����r|ن�]f�^��4�ʓ ���, �ӂ�5��f��-�w�г�����.�\4,a��0^��Ձ3��H����ƙ����5s��}��*�xU���A��3/�!��͆E�����򘎽���l�Q��,���U2U��ߜƃD.���5��m�r�2��FL1�����_�����q���u=�D!{К�@l,���~lf���2
��}���̯A��|�dG�}�/h����� �$/�X,�Y-���$���A�]��HW�"�xP���j�,����J�l��K�	C�m!ͅ6L��|'9��������}�'$���5aJq+�-��6UV� �0�u�.ˆ�¹����a�,�KLZw��r����0H�<A��Fp��jX��_F����`yl����Q���"~s�X����>�A�� ®�	3~����,-����6�ǅw�t|QcZ'�i+�V-���XP��X��*E=��^�
�4�Zf|�8� 1���.͙e��V u,��3��'v	� �t9q{���O�M2���h�oc�ݻ���)XT$#�ؑ�ә�4|K]���C1��o/;�#�[n.Ҷ��~�2Ar9G�>usH
�L���w�����l���v���6��.i��U;�d}*��G�- WH�'���m��F�t|ٟA,��p�~���$��m��~E�d.�`n7MI�WEd9���m�@R�����߫��I�	|�m�](nY(iy�{��[��g|f)��O��p J]儳��s!ރE%�s��;��Etht):�d���q�)�'��7C�e��NX����t�*����EM��t��x*]7�}�@4�%W���_�65ǉm��tk'��sm9���"���4�$�¥gf���5m��l���.�M>ݭ�NH���B�B�c򍵪{;�/B�v��>:��䐤B�ٯ�FTf�z1{��N�}#_��퇧}-�P:0�߹H�*��Ή{%����H���GD>A"�����h�j�&Z�����zZ�W.@YS-�o[>
���X��������~���xt��>-h������{�LY}���ʬ�8����7�D��iأ(._�ս�_ZMٻ��� /��
F٥��]�����4��:�|��m	GȜ&������<�Q�r0l�}����,�\X��OiKl�X8�9��u�Х�Id�5�����D!%h���]��r��Aޮ�A)��!᫜�fȝ��L�an�b���}b
�$Q Űd����)3"v�2Go�V��H=��a�24�5G{�R]D+���P��:���!~v���jjd��ym�O�}���hA)��x��5*����ʛk�v#)	[ý>�����U�ɽ�٤��ɾ�[-�Z�(�[��+$��袽/�������w�qE`� �6�a�!��ot�NQ�?�)4��۔?2�� m�g�RL�vpdY�
3\��E�kI�@��	F�\8B���dX�[\��+�О��ڽ,ki ����=H�1ƀ�q�1��(����^p#������2aa9����L%�)`�c�W���b
��!��u'ziII�'�6�F��Њ� �Aa�֜MB`O���m�zȢ܎jm)�C�<+qn�)x��mݱ��pu���bq����'圩M���b�)�[cKm!WY��)��G�׼>�7��D��nQ�Mޗ�X��2�"�%�����5�-zU�T�b6�Pq@�dY��H?�%��s��L�[PiT�5���zH�(���˨����Zm�"t]E����p7F#9_�"���O��"l�o�����:Ep�g��~k\X�G�ܩ�����哭'�l[���?y�w47�P�ޜ�����.�O%�(.T����,�$�:�?ݏ�yh���.�͌l7��i*8��VX�S�{f���3��Q(Ҷ̌��򟅽gA��50�։����Qt�b����t��ef��+E!6��~H-F$�~�0s%���0��#?yc"&2 �z7U5�;�5k�l7�X�������]��c�ُ�c�����͂8=��0^�R���yE7~SV.I�1OC�����w�y%?,�KI6�ۉt��;���
� ���+�RF=vJ?93{�4�-Q�)jk�˰s�.�����b�4o5f�ࢹu	�!5��>F���ܦ:�����졍��5�`�켍7�Q�`��8����&����9択�fߍ\�J��s��9�ـB��6��J֭��PϭZ��dh�ԭ��^b�2���Q|�B/�ô_Xj�G8�w�E���M�N��R��+�O!0Z�t�@�m\��Xv]q��}���2��nu��un��%���.9��"`�5�%�1"W�+D���[	�%q��v��@lײcΤc�y�	1A.��>��Cw�ܲE���]{��M8�v���:�M+����â�UԖ	�]H�VqrT����r��C��z2ѽ�앧�����u�^�q��-|g�� ���:)*�פ��Y�>��M�%���&o?���ΣMM�!�L���W`�v�UD����[��capnJ��ˋ
�Ѽ3N��18<q�Xf�.62�z��7��c?��˰��Y���%9�m�f���% o|�� MD4Jz��,�V��L���c�.�%�����u`�}�d̏5����=��r�:�K�3יLÄ����x�>�fZڇ5��ւ�0�S�I+b�u1#H��6�����j4rX�f�x9
 y
���q.)�P���3]��t��)�2�x�d���ݓteY��0SLHXoE�j
vnJŵw��?RX���!����                                                                                                                                        ₆H          (  �    �   X �    ₆H      
 1u  �  �2u  �  �3u  �  �4u    �5u  ( �6u  P �7u  x �8u  � �9u  � �:u  � �    ₆H           �   �" H  �          ₆H           �   �( �  �          ₆H           �   �+   �          ₆H             �, �,  �          ₆H           @  �Y �  �          ₆H           h  (i �  �          ₆H           �  �q �  �          ₆H           �  pw 4'  �          ₆H           �  �� 4  �          ₆H             � �  �          ₆H          0 �    ₆H           H  е �   �          ₆H          p �    ₆H       	  �  h� �  �      (   /   ^         �                       �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                                                                                                                 83333333333333333333333 ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� ?���������������������� 8������������333333333  ?�����������            �����������             ?���������              ���������               ?�������                �������                 3333330                                      ������  ������  ������  ������  ������  ������  ������                                                                                                                                                                                                                                                                  ?��  �  ��  �  ���  � ���  � ���  � ���  � ���  ������  (      >         l                       �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                 s33333333333333 �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� �������������� x�������wwwwwwp �������         �����p         �����           wwwwp                         �����������������                                                                                     � ���������������    (               �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                         xwwwwwp �����p �����p �����p �����p �����p �����p �����p {���wwp ���     wwp            ��  ��  �                             ��  ��  ��      (   `   �                                      �   �� �   � � ��  ��� ��� �ʦ       """ ))) UUU MMM BBB 999 �|� PP� � � ��� ��� ��� ���   3   f   �   �  3   33  3f  3�  3�  3�  f   f3  ff  f�  f�  f�  �   �3  �f  ��  ��  ��  �   �3  �f  ̙  ��  ��  �f  ��  �� 3   3 3 3 f 3 � 3 � 3 � 33  333 33f 33� 33� 33� 3f  3f3 3ff 3f� 3f� 3f� 3�  3�3 3�f 3�� 3�� 3�� 3�  3�3 3�f 3̙ 3�� 3�� 3�3 3�f 3�� 3�� 3�� f   f 3 f f f � f � f � f3  f33 f3f f3� f3� f3� ff  ff3 fff ff� ff� f�  f�3 f�f f�� f�� f�� f�  f�3 f̙ f�� f�� f�  f�3 f�� f�� � � � � ��  �3� � � � � �   �33 � f �3� � � �f  �f3 �3f �f� �f� �3� ��3 ��f ��� ��� ��� ��  ��3 f�f �̙ ��� ��� ��  ��3 ��f ��� ��� ��� �   � 3 � f � � � � �3  �33 �3f �3� �3� �3� �f  �f3 �ff �f� �f� �f� ̙  ̙3 ̙f ̙� ̙� ̙� ��  ��3 ��f �̙ ��� ��� ��  ��3 ��f ��� ��� ��� � 3 � f � � �3  �33 �3f �3� �3� �3� �f  �f3 �ff �f� �f� �f� ��  ��3 ��f ��� ��� ��� ��  ��3 ��f �̙ ��� ��� ��3 ��f ��� ��� ff� f�f f�� �ff �f� ��f ! � ___ www ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���   �  �   �� �   � � ��  ���                                                                                                                                                                                                       ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��������������������������������������������������������������������������������������������  ��������������������������������������    �                                                                                                                                                                                                                                                                                                                                                                                                                                               �������������������������          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �    ��������   ��������   ��������   �������������������������������(   1   b         |                     ��� ��� h�� P�� ��  �� 8�� @�� @�� X�� x�� ��� ��� ��� ��� ��� ��� �� ��� ��� ��� ��� ��� ��� ��� P�� `�� `�� p�� @��  ��  �� `�� ��� ��� ��� ��� h�� P�� p�� X�� 0�� P�� h�� ��� ��� ��� ��� ��� 0�� ��� ��� ��� @�� `�� ��� ��� ��� ��� ��� ��� ��� h�� �� H�� p�� ��� ��� ��� p�� X�� @�� 0�� ��  �� @�� @�� p�� H�� p�� ��� ��� H��  �� 8�� H�� p�� ��� ��� ��� ��� ��� ��� 8�� Hx� p�� (�� P�� h�� x�� ��� ��� ��� ��� ��� ��� ��� Hp� x�� `�� ��� x�� �� Xhh ��� ��� P�� ��� ��� �� ``` ��� x�� `�� H�� (��  �� h��  �� hhh ��� ��� P�� 8�� P�� X�� ��� ��� ��� ��� (�� phh ��� @�� p�� ��� h�� 0x� ��� ��� �� ��� ��� @x� ��� 0�� @p� Xpx @�� ��� Phx p�� ��� ��� `hh X�� p�� ��� �� ��� h�� x�� ��� h�� �pp H�� @�� `�� ��� `�� P�� 8x� 8�� (�� X�� 0��  �� ��� X�� (�� 0�� ��� P�� Php x�� ��� x�� H�� �� ``h H�� �� x�� ��� H�� ��� p��  �� ��� h�� P�� 0�� �xp 0�� ��� ��� x�� `�� X�� 8�� �� �� `�� H�� �� �� @x� Px� hpp xhh  �� ��� X�� @�� 0�� �� 0�� hh` �ph (�� 0x� `pp ��� �� Pp� X��  �� (�� �ph Xhp (�� ��� l�� T�� ��                                                                                                                                                                                                                                                                                                                                 ����                                               ���䥂��                                           ����q��_���                                     �諹���qԚ�����                                 ��٧��ڴ��U�q�������                             �i�������ϫڹӐ��������                         �i�����������������U���_�����                    �i���������������������U�������                  2 �������������������������Ӑ��_�                    �Ąń���������������������������                    �γ��������������������������ꁎ                 K �έ����������������������������                 úJ�έ���������������������������q�                 B����zttttttttttttttttttttttttt���                 B����zttttttttttttttttttttttttt��*_                 B�a��>tzzzzzzzzzzzzzzzzzzzzzzzz��M�                Bu���%4444444444444444444444444t����                B��c<$4444444444444444444444444t�cԯ                B���:$%%%%%%%%%%%%%%%%%%%%%%%%%t����                B����#%%%%%%%%%%%%%%%%%%%%%%%%%tp��                B��L�#%$$$$$$$$$$$$$$$$$$$$$$$$z�sq�                B��V:=#########################>�<�                �e�U5=========================��;	_�               �e�KeCC""""""""""""""""""s����               e�HUWe�Q5�vvCswC���               fs�GIa�b�W�YZv<�vX��               \s444t�?�HIa�c5vCCCCCCCCCCCCC;�Y��               �5=%4%%%%%%%4mI�\hvvvvvvvvo�h0q�                :=%%%%%%%%%%$mI�Q�vghggggggow�q�                5"%%%%%%%%%%%$`ܜ�W�Y�05�ghvil               QC$%%%%%%%%%%#"$R`GSIa�b��Q5�5D	_               �"%%%%%%%%%#Cooo"""=$R`GS�JL�OP                *ZC$%%%%%%%$C5,	!�38/5;;"==#%?@'��                 �,###$$$$v,'( ��+�./5�B                    �f]Cg�       �B�                        �M!8O                                         ��������                                                                                                                                                                                                                                                                                                                                                        ������� ������� ������� ������� ������� ������� ������ � ����� � ���� �  ?��� �  ��� �   ?�� �   �� �    � �    � �    � �    � �    � �    � �    � �    � �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    � �    � �    � �    � �    � �    � �    � �    � �    � �    � �    ?� �   �� � ��� � ���� ������ ������� ������� ������� ������� ������� �������     (      >         \                     ��� ��� d�� ��� ��� ��� ��� d�� x�� ��� ��� ��� ��� ��� ��� Lx�  �� p�� ��� ��� |�� P�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� d�� 8�� <�� ��� ��� ��� ��� ��� ��� p�� X�� @�� @�� 4�� L�� x�� ��� ��� d�� ��� ��� ��� H�� 0�� P�� l�� ��� ��� ��� ��� ��� ��� ��� ��� 8�� ��� ��� ��� ��� t�� p�� @�� P�� ��� ��� ��� ��� ��� ��� ��� ��� ��� D|� ��� ��� d�� X�� \�� \�� P�� L�� d�� ��� ��� ��� ��� x�� Lt� d�� t�� 8�� d�� t�� ��� ��� ��� ��� ��� ��� ��� ��� P�� Tlt `�� ��� ��� ��� ��� <�� Xhl \�� l�� ��� ��� ��� ��� (�� Tdh L�� X�� ��� |�� ��� (�� $�� @�� ��� ��� |�� 0�� ``` D�� <�� ��� ��� ��� `�� <�� Dp| x�� ��� ��� ��� ��� H�� D|� 0x�  �� ��� ��� 0�� Pp| 0|� d�� $�� ��� x�� ��� ��� |�� |�� �� Thp lXP `�� <�� ��� x�� |�� |�� ��� ��� �� Thl d�� ��� t�� x�� ��� ��� T�� 8��  �� �� \dh 4�� ��� l�� t�� ��� h�� L�� 0��  �� (�� 8�� @x� Dlx Xhp ddd h�� L�� ��� l�� x�� \�� D�� $�� �� (�� 8�� Ht� Lhp Tdl \dd l�� d�� ��� T�� 8�� $�� �� (�� 8�� Hp| Phl Xdh `dd h�� $��  �� �� (�� <|� Llx \lp                                                                                                                                      �ځ�                           ���������                       ���������*綁�                  �c����������k���              ��i�����Ŵ��������\���          �3�Ľ����������~������          �3��������������������          ܮ�������������������z�         �������������������ԫ�         ��������������������ӥ�         ����MMMMMMMMMMMMMMM��*�         ���,����         ���,,,,,,,,,,,,,,,=�i��         ��r,��<<<<<<<<<<<�h��         {{K-vu||t}}}}}}}t~��         lmnepKr
-twxyz         ]^_`abcefg----Wixjk         K<==�OOQRS
TUgWV�Z[\         "<,,==>?RADEGHIJ         +=,,,-./01233n6789:          !"#$%&'()*           	
    �c                                                                                                                                                                 ����������������������� ?�� ��  >�  >�  >�  �  �  �  �  �  �  �  �  �  �  �  �  �  >����������������������    (      "         �                     ��� 2�� 0�� .�� -�� 5�� ��� ��� ��� ��� e�� �� C�� ��� ��� ��� ��� ��� ��� h�� �� �� � }� |� |� @�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� v� Nl{ 9�� ~�� ��� S�� F�� H�� D�� a�� w�� u�� s�� p�� X�� x� 0r� 7v� 7�� u�� U�� ��� ��� ��� ��� ��� ��� ��� ��� ��� b�� ��� x� @q� 4�� j�� 6�� ��� ��� ��� ��� ��� ��� p� bef 1�� b�� :�� ��� ��� ��� ��� ��� ��� e�� ��� o� `fi ]�� 7�� ��� ��� ��� ��� ��� |�� _�� ��� m� `fh ,�� ^�� ��� ��� ��� ��� ��� r�� X�� ��� k� `fg *�� ��� w�� x�� y�� i�� R�� ��� j� _fh %�� P�� %�� m�� f�� [�� [�� Z�� Z�� Y�� L�� <�� l�� i� afg %}� $|� "z�  x� u� t� q� o� m� k� i� h� f� f� cfg eff cfh bfg � � �3  �33 �3f �3� �3� �3� �f  �f3 �ff �f� �f� �f� ̙  ̙3 ̙f ̙� ̙� ̙� ��  ��3 ��f �̙ ��� ��� ��  ��3 ��f ��� ��� ��� � 3 � f � � �3  �33 �3f �3� �3� �3� �f  �f3 �ff �f� �f� �f� ��  ��3 ��f ��� ��� ��� ��  ��3 ��f �̙ ��� ��� ��3 ��f ��� ��� ff� f�f f�� �ff �f� ��f ! � ___ www ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���   �  �   �� �   � � ��  ���                       ��������������     ����������������   �����������������   zo{t|}}}}}~����   nopqrssssstuvwxy   bcdefggggghijklm   UVWXYZ[[[[[\]^_`a   JKLMNOOOOOONPQRST   :;<=>??@ABCDEFGHI   *+,-./0123456789     !"#$%&'()            	
                                                                   ��� � � �                                 �  �  � ��� ��� ��� ��� (   1   b          '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��  
<hl [C   .                                                                                                                                                                 �� ��i ��� s�� Yv�8K�� �t   `J   4   $                                                                                                                                             �� ��y���N���,��������� v�� _�CZ�%��zgQ   :   (                                                                                                                             �� ���&�������j���Z���T���C���-��������� y�� e�� Le� (6�
�  � mW   @   -                                                                                                            �� �¥(�������x���m���m���h���c���^���Z���J���5������
��� ��� q�� Uq� 4F� �  �  s   ]  G2   "                                                                                         �� �Ĭ)�������}���o���p���p���q���q���q���m���g���a���\���P���<���&��������� v�� [z� >T� '��  w  b  L7   '         
                                                                �� �ī�����������r���s���s���s���s���s���s���s���t���t���q���k���d���_���V���C���0��������� y�� c�� H`� *8��  {  h   T   @   )                                                           �� �«�����������u���v���v���v���v���v���v���v���v���v���v���v���w���w���v���p���i���c���Z���L���7���$������ {�� i�� Qm� ;O�  �  p   <                                                        �� ��� �����������x���y���y���y���y���y���y���y���y���y���y���y���y���y���y���y���z���z���z���u���n���g���^���R���>���+������x��D\�   ^                                                        �� ��� �����������}���{���|���|���|���|���|���|���|���|���|���|���|���|���|���|���|���|���|���|���}���}���~���{���r���k���Y���+��� e��  m                                                        �� ��� ���������������~����������������������������������������������������������������������������t���;��� m��  x                                                       |�����������������������������������������������������������������������������������������������������������������������z���G��� |��  �   '                                                �� FY%����������������������������������������������������������������������������������������������������������������������~���N��� ����3                                                �� g�-%���'�����������������������������������������������������������������������������������������������������������������������T������ "-� @                                                �� ��B%���'���u�������������������������������������������������������������������������������������������������������������������W���"��� :L�  M                                                ����A*���-���c�������������������������������������������������������������������������������������������������������������������^���9��� Jb�  Y                                                �� ��BB���F���d�������������������������������������������������������������������������������������������������������������������d���O��� Xv�   d                                                ����KR���W���i�������������������������������������������������������������������������������������������������������������������j���d��� e��  p                                                ����hQ���W���X�������������������������������������������������������������������������������������������������������������������q���y��� q��{   !                                             ����|Q���^���B�������������������������������������������������������������������������������������������������������������������x������� }��  �   )                                            ����{c���q���@�������������������������������������������������������������������������������������������������������������������}�����������5                                            ����{}������D�������������������������������������������������������������������������������������������������������������������~���������� #/�C                                            ������������3�������������������������������������������������������������������������������������������������������������������~�������5��� ;P�   P                                            ���ª����������������������������������������������������������������������������������������������������������������������������������L��� Mh�[                                           ���İ��������A���:���m�������������������������������������������������������������������������������������������������������������������d��� Yx�   g                                           ���İ������������U���1���,���?���Q���[���n�����������������������������������������������������������������������������������������������}��� i��s                                            ���ð������������������������}���f���P���B���/���(���9���h����������������������������������������������������������������������������������� t���   #                                        �����������������������������������������������������u���2���T������������������������������������������������������������������������������� ���  �   .                                        ��������������������������������������������������������w���+���b�������������������������������������������������������������������������������<   
                                     �������������������������������������������������������������r���6���1���V���k���{��������������������������������������������������������������6H�D                                        ����Ͷ�������������������������������������������������������������������u���]���K���4������'���<���O���r�����������������������������������3���Ha�9   
                                     ����sj�����������������������������������������������������������������������������������������������v���_���I���6������$���B���A���k���u���!��� c�u                                           ��  ����ΰ���������������������������������������������������\���5���[���q��܈���������������������������������������������j��� ��� \z� ��� ��p :O                                                ��  ��uX�����������������������������������������������^���d�� :Q= 9M0 ��I ��c ��� �â�ɷ%���H���f���z������������������������  ?    ��                                                      ��  ����Τ���������������������������������������}���x�� ->G        ��  ��  ��  ��  ��  �� ��" ��? ��[ ��y �× �ƭ ��� ��� ��o                                                                       ��q���4���R���m���{���������������������,��� Wxg                                               ��  ��  ��  ��  ��  ��                                                                                  ��- ��: ��[ ��p ��� �ġ �Ű ��� ��� �g +9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ������� ������� ������� ������� ������� ������ ������ � ���� �  ���� �  ��� �   ��� �   �� �   �� �    �� �    �� �    �� �    �� �    �� �    �� �    �� �    � �    � �    � �    � �    � �    � �    � �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    ?� �    � �  �� � ��� � ���� ������ ������� ������� ������� ������� ������� ������� �������     (   !   B                                                                                                                                                                                          
                                                                                                                       	4   3   &         	                                                                                                ��  m�$^~l"-�	�~jS   <   )                                                                                        �� ��U%������~�� f��Le�(5�
��oY   B   .                                                                         �� ��sK���i���_���J���5���#������ o�� Vs� 6G� �  �v   `I2   "         	                                            �� ��wK���z���t���k���g���c���^���R���A���-������{�� \|� @V� "�  �  x  e  O:   )                                      �� ��w1������z���s���t���t���t���r���m���h���a���W���J���6������	��� d�� Ib� *9��  }  c   9                                �� ��y*����������w���x���x���x���x���y���y���z���x���s���m���e���_���U���?���(������ h��BW�c                               �� ���+����������{���|���|���|���|���|���|���|���|���|���}���}���}���{���r���i���_���A��� h��{   !                             �� �ì#������������������������������������������������������������������������������_������  �   *                           ���ͫ�������������������������������������������������������������������������������`������	�5                           2��1�Ӭ�������������������������������������������������������������������������������g���+��� %1�A                           1��/�Ӳ(�������������������������������������������������������������������������������m���9��� 6G�   N                           ,��+���)�������������������������������������������������������������������������������v���Q��� H`�[                          7��6���0�������������������������������������������������������������������������������|���d��� Zy�   h                          G��P���J�����������������������������������������������������������������������������������|��� g��t                        w� ?��_���^���������������������������������������������������������������������������������������w���   $                    u� [q`���a�������������������������������������������������������������������������������������������   ,                    ����2`���s���[�����������������������������������������������������������������������������������5���� 8                    ����Bu������^���G���J���e���s���|���������������������������������������������������������������L���%1�D                    ��	��B�������������������}���g���V���C���C�������������������������������������������������������k��� 9K� P                    ��	��A�����������������������������������h���P�������������������������������������������������������Kd�X                   �� 
��7�������������������������������������������S���R���b���o���������������������������������������c�� J                    �� ��a�����������������������������������������������������������}���d���Y���H���E���\���e���f���f��� z�� #                       �� ��s�����������������������������������X���<�ƫ^�ܹz��̓��ӫ��ܷ������������������B��� d�� u�q k�,                        �� ��O��ǹ���������������������������\��� JbW   a��  �� ��# ��E ��d
��~/�ϣM�׵W���F�հ Xw1                                            ��[4�К@���d���w��ڍ������h�����f                                      X��                                                                     ����1��> |�$ Pj	                                                                                                                         ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����   �����   �����   ����   ����   � ��   � ��   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   ��?�   ����   �����   �����   �����   �����   �����       (      "          �                           !   -   /   /   /   /   /   /   /   /   /   /   -   #   	5	o	����
�
�
�
�
�
�
��q   8=V4{��w��s��q��n��l��i��
g��e��c��a��_�� ^�� T}��w$���P���&���m���f���[���\���[���[���Z���Z���Z���M���=���j���W~�
�*���^���-�����������w���x���x���x���x���x���y���i���R�������e���,���^���2���������������������������������������r���X�������f���.���]���7���������������������������������������|���_�������h���1���b���:�������������������������������������������e�������	j���4���j���6���������������������������������������������������l���7���u���U�������������������������������������������c�������v��#Z9���~�������S���F���H���D���a���w���u���s���p���W���u��`��s��"0@���������������������������������������������������p��   N       C���������������������������j�����������}��|��y��        2��5�̼����������������e���e�u���� �� �� � y�             3�� 3��2�˾2���0���.���%w�c                                          3�� 2��2��0��.��%w�                                                                                                            ��� � � �                                 �  �  � ��� ��� ��� ���    
 //   H  1u   �  2u     3u``    �,  4u11    �  5u    �  6u    �  7u11     4'  8u!!     4  9u     �  :u      �4   V S _ V E R S I O N _ I N F O     ���                                           D     V a r F i l e I n f o     $    T r a n s l a t i o n     	�4   S t r i n g F i l e I n f o      0 4 0 9 0 4 B 0   4   P r o d u c t N a m e     F U C K   Y O U     , 
  F i l e V e r s i o n     1 . 0 0     0 
  P r o d u c t V e r s i o n   1 . 0 0     , 
  I n t e r n a l N a m e   t a s k     <   O r i g i n a l F i l e n a m e   t a s k . e x e         �� �� �� ��     @�     ����|� @�                     kernel32.dll      LoadLibraryA    GetProcAddress      VirtualAlloc    VirtualFree  ��p�t���s��v��r� ��6� ]|$nWخ  �H�0�
U��r�u4<E9H�8e�g� 3�BSV�pWA���0�}y��E�ȸæh��?KOu�6��E>]��}��U�@���t2�W���7��>j�y���Y�u~`U�6����7*Id�u�9M;w�3�_^[����r�#��M��V����
�<�=��s$ȀM�0:�ʺ�應"9�>�����9u<���p���+��0S�7(hu���#��jY*M�����F�
�B�i��� }����l�zl��@�|+P�Ƅ1,��e��u��эgd�"ؔ�@]u��@��@u	��s��:�؁҉1��͂���)H+Ƌw`Μ؉�T>tg(��x��s��ap ��u�6D�>s*b���n(�k�g2|�����$�U�<�	+A�#23
m���<�������꒜�[ŴT�ύ&��CH��F
�C�3�j�2N��0Hx72�}���(�E���	���"������
6W���0U�VVQ����94��j�[��������B��ǦP4��6�S���&��X�UC�sGDU�SH,�D����,�Q?BUH{3ɤ����L	�~�6�T����;�[)Ę+q *�p�"�`�&�T�x2�HzT퐺�����UI��uY��b�vkQK<I���$j������n#��U#��%S�&
\�$1m3�cN�!��eE�։�`���a&�q\4f�(���e)�b���AE�&_���]S��"�G��;�����G�C�ɉ4���G�|l�.\�6�������cP�>��+����,"n�z�og��mF��rjxY�(�X��9��inI����]��"ҵ9�h�H� u���@���p��������&��,¾�}X��a@p��
��C��~;���9�qr)�
��uЍ���L
���"�gG�2}�O���M��ڹ����r�B��Jf���n	�|?�R }�C��&����Tq�;�w5!`�+�ϊJ�D>FA��	A���Jt;Qr庠�9���w��3�@ÚK"�p�(u� FW�j	Y�u�<_|phKZ������}}����B�ä'
�� ��H�Pj�Wa��8��~?>S�ʃ6�	�}�7�~���QK�P_^��8�UH�P-XpT@,g(
P@���D�XF%$�5��Dh4��$���|�aA6���6�@�"�=��!S.WVP ]��LT��C�F���+�޵V�v����/b2�����	{Ht �sD���4�#��S{@���w��X/�o1���Q�F���0�N,��+Kj@�s�QF'�7!��'V�U�߈r���6���(@�U�ɐ=��4���#����Q�FG0nt{������*Du�D:�-��W�t�R'��CQ��f1P"?��LB&B���A�R�?Ұ���bj����fH1��7$�%Du	C��K@��������4��%¤��(�W�7�(<��3�;�@F�]	^_[Ð�����p�[��?�`�Q�H���T��X(~�r�L��vtR�~��P!��3�E�Z���L�a�uŚ�����Т͉�f`��JI�������L��t�VC��\5>��X<t
�H�0	P�:.����F��u}�-�I���zkl>�@>^ 6u�;�}y4.F\ �U�,���}t�Ȋ�u*:f����&����/,���`A��^Y��Ft5;*�0��B�)��x^�Q��9�!4`�fvR���Y�XI?&W棳��XA���S'rPޅ�C�!HtM��s^}(KY�8����-�����{����R��>�!�	�Zi';�2=i2��u����E��G��QRVF��#�"֡��L�}\�&jnH+�
6�TL^ �b|X	��1�H�RdK�K���/�Q������@t�%��F�)�?6������Z���;}u��Q��O@���H�9��+�I\q^�'�"�@�-I-@g��F��)�h"I�&9\(��t$�DC�QN�h�~3��!{�PWQS��ǂHF���@��N�p�msvrb�2���E�K�[��!��F"���XN�[9�҃OӑY��p0N���Nc����2�}��U����������Pn��?a�tDRH��%B	%r#pj-��A��f��Q@�YI�4Zh�loXM�rKTE�����\���*o���*0+�i��H;$MfA��}60k��m�� �b@<��H�|��'���X�`9�Q�vPi���:� ����,��Y�(�rǥ!ed�VR�z"ȧeH%3S�.�!�4J�{ �����-���
V4��ޙH]�Ap�lic:aton er�n|)�� �u��.The��<vcd�%s5�l��n�t�b_va6�i�d�SDL�BG5f�d,7al z3W�*WN'c��,us�32M�y=ag�BoxAw��1xtf�k8�6l?ExitP&�L�C��hHa<nd~�Ozp�XG�tzM��lM�|Virt��A�c�7�v�2�	�$�J���fm9�	D�P�<H�0z4I��	���wl `�t$$�|$(���3ۤ��m   s�3��d   s3��[   s#�A��O   �s�u?����M   +�u�B   �(���tM���H����,   = }  s
��s��wAA��ųV��+��^��u�F��3�A�����������r��+|$(�|$a� ��   	  �� H� L�   @ @� D� �	�C���� �A�T$�R���+ʉJ�3�øxV4d�    ��USQWVR��W �SR��j@h   �sj �Kʋ��Z��PR�3�C �K �C�K�KʍCPWV��ZXC��R���F���+��V�K�N�׉�? ���KZ��h �  j W���Z^_Y[]��                                                                                                                                                                                        