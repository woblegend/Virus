MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                                               PE  L n��G        �   P   .      �1      `    @                      �     ��                                ��  <    �              �  �                                                             4                          .text   �O      6                   �.data   �*   `      :              @  �.rsrc    `   �   `   B              @  �                                                                                                                                                                                                                                                                                                                                                                                                                                        ��=��<}9�rm�(JnQ����-���zh�5�Im��c�����i�Bۏ�G>3����L�q�uG�6)�g��_L�FfD=պŵ`2g:��"��-[���H�X^��7��<B�v�єT����69>�SJ0������Ί���h�^�����O��"���Vb~�O�N牅�#�+q��XZ�?��|kz�-;&݇'z��=r���[�3s d�R�L����}Jqz�S��Af�l#�>���`ڿ���3�Y���K<�}I��w������S���뺇�#���>�~�~�]���� �j�d̓RK�[ƄI��u����z�q���0IiC`� i��O���ݦ�ZM���z,�=��}�k�� ���pYR�����	�>�.�p5?%�B�m��ϥ���b.[_,�H������_L�����R���@ɴ��)��*`ALw�3�	����2�Ŵ�M'&)%�=dQt�pצ��'�k�o�\��P���(	�q�NI���D�F����ǙOTlBn��ا�*�l#=Ы��� h�"nĵ'Ƹ�g��v ��G��0.��5}��`��ʳ['r��mSZSy��mА	fX}���h��.dC�,Q哘&�Hִ|��O\�%-h`M/����� �;KK+��O�<k'Z~�j7����8�Ǿl#4�Yd�?��:n�Le��-K;�~>o�Ӫht0;S$�I�T'~�$e$��^�u���DE�<8�%1*�~H6�Rj����i	�c?����e��f
�E��t����)�=/ì�ٔ���wy��kO�}8Ƃ��o�k�D���&��e��,��"�m�06�]:��+�Y@��h�<%������-��W�ϓ�;�E:P1�r)w�W���[��\=����*~o�_sb��w5!,�/�� 1�#o������̠����������)m@LJU	�p���7D
(����ڠ��8i���r<��v��T���.��4�;��Jd�8V��~�$������"%�k�z��c��	�s�qg��DT�p,�0�f��7�5���N��p�&��@N��E�,���HՇ�H�+�����_���Z����5m2z�:��a���4�j��MZ�Fd0(-g�o�u8al����c8V)U����.���L"�/�OC?���M_%<�p�J�A����DY2f�L"_�g1�)��@���^e¤��Z�E�� D�ۀ�^1�:��J��+�hN2<s+��eH9S%E�̢�hG,�=l5�_�}��M�F;P��u7�\F�7+��,�{���NMW
�KM�L���$� �=���?�|���F�����B/��j���,  n��w7�C�����
��;a�Tc���et�/@襹E)�a����D��>�M��f$Sj�TA{}	*7ȲUx�ՌL�p6���9V���b��n�z� ,��:�
^/�����.�����l�f��ŷ�x/ƣ�a�R(P�Q�7[�p�y�����/}�\�<�~*b���w�&�E��^��ݖ*Zd���;}�{
o�um�N����x���+�d�D�ח��7�Tz���y���pfKz��8��S"#�L���N	��
��n�=���� g"�ЯkޠD&^�Ba��&�'������x�{�Y<�o!��2^��6?	q�RzN��FO����gY5^�+\�]��W�� n����>�D.`n	q�8��H��k`3#��%ވ��5�'�Ϫ܅v�e� �s�bJ	�j�c�A��.
iPB�{���;NpOx'��<�]����f�n�K��.�e�����O3v����G�!�
�1�J)S��'t"6��]b ����%�'��g�8��v�Rf��`[y���f��!��b���2�MV�g΅��-��M��1��g��P��򟹳XmRA��neXaͭ��+�Z�blj�qi����~��8x��.�D\�,�0נ�,M�=4�ۡBUى�A%�LW�c闃M�Tl��iW����3R����x0��^�����Qs�/l�!��I�d�$I�C�<�����2�݂�ѱ�4��j�����h�ָ Ls�\�99N��R^�=��z,I*�p@�(��9���A�`���[���wL����Ki��3IGu�� �H��˦HW���$"J̛�j��� Õ�O,H��_"岂l�Q|%�C���ͺ�Ep�#� ��@.k�XX�p��sc�E�X���qi��a���ć��#�]St���t��E��[�� ��]�'��S�h2t��0�A����?h�:�`B+k4�l��]>�w�ʠ͌�?6�]>`���:�9r�Sp|'B����������8g6W��� �C!��8�_םl]�_[��TJY���=���&\-�S�"3�J�;�����m={�V���H	^ɇ�>q�Qj��҇�䗷�=*g6b��]=�䔫7#ԗ�K=v 1�M��5iJ+�F�"�9BQmG�`�z�����[���$ <�Kے姧�-���l(��Q���1?���QI�5W�K�Q�Vʡ����~�������e݄�)}��!��7��
e�,�[mwS��RZ�KY�?��G�h��''kA�^�B�*lα��v��E�#xr��T�v���(�/5�6w�8�`Q5��Ƿ�A�⼝W�2 a�����]�+J��Hϖ�CZ��_�7�}��|��/���ZE�T��k�]�t[1n�M݈�Ѡ�ـ�_t���K�hʩ]�z��l\�y΄[6&\��4d�>�=�;/o��
%9L��Η��u��_$L?v�o0Ei�(�|J�G��װ�4������u�(��:6׾<%��Pg蒵�q#�]%Ѕ��X�詓흉ԉJ��t���LLK�L�ѽ˄���Ek��>�v�W}-�w<�b_��ѩ	o=u�G�􊨌LG�X ���d���şq�dd!����m��N`�D�1�hOP�G��ovx�ҽ��yN��Wu��?p�#qU�\��F�qn����]����4$�՝��	3� �,��|�4�Č��d��fE� *�s�`�U�"�T�ݍ���jm�U$v�˂���c�����C������f�^w�(���y)@�ٍ�(��`�ϛ�p�q����!��>C	0|[g1�w�TX�1~�3�K�x��^ĕ�r�w��A����\�T�MqF�����0G���g��fe��� �_� �O,�N��/��� ��͎[�r�_�C���B�xk2���6���q!�v*����rj-V����2�dJ��%B��7@Í���Fg$܆
��!|H&Zj��/�D���5���pn�b�A�x�Wǡ��CN��Cs��.i�y&�f#A%n+����x�\/��`��:[�/9p9�H�r;*
��	�=��j��>`;\A�!A��=�Wa��8E�:,���l���:�W��(����H�4�� 2Y�P�lx��i_g�I#�f$��k�����WM�uEǘ�q��yn����C����gmE�v��Gi���G�/������
��:�?J��W0������r�x[X�w��$u�H��X��3�;O�LԑE�Y:��?�n�᚟����47*�.1F����vXB�����pi�2�����J�7	���M��gJ�������2ɺuD0oi/���&Өξ˄	Qၯ��1�aG��ڣc����]�`J��W	]�r��3W��n>R�|��h7�S���ɡu�b>J��9��lm�<;w���M�jP�LT^�<ƭ�>�c�1��C&�{p!���K��h��t18���HN�L�SC�C*�/��J	��3����dA�w�-�b��@0�p՟4B���-���U�V��L�5��HR��
������eZ��)�n�g"�Bo����Ԇ��t�f�>s�F�&]�!��G����o���ru���@��"��������j]��7v�y�^e��r�m7��>#3��-U~��{D�\��
��f�أ�>:w���6�aZ�`đ�ۏP|Kl�Dc��n�Drx~M�W�w��>uJht�����}
u.I�ڤuR�����f�� 	5�ݒ�V@����F�;��<�z�_ �֯�xK���nn�&W�65f�
��IxT��|*XdF�(l�hy�wv�#r:�QeihK]F����yYW�o�*���=V	^�?�u6�Jn15Ѿ�-Z�����"� �9鏰�!�!|y��� ��A��Kw8�S��	D�v��"���)��¨)�)��;�Ԏ��z�(����[(�i�!�	���A'q�kQ��#��覧!~RU�ׁ���joS{�Ҳ����F��Xq�������2��PG����nq��2���:�O�c>xT%w� �s� ^=L�`��K[�\2�Ɏώ��FФ�Uͤ���E�{Rr
%��ZM�hC���w�V����R6J�ގ._�1@!Ȥҏ!�ȋ��/�7���HH��\���n�q���IG7�4ǎ�PM��-����^"��n�#y��MY�$�T{��H�񖽋K��0 �����z&����N�|��B^��Eg���}�e8-�[�(Z�l��T�GD���P��?ܬB][�<Aj��TA�������"�����[�JM�������|ӡ���FjI�z�|��OI�ؑ[ժ2Y�4QX(ŧ��ꇂQ;NBx���rx�e�l��S�5�o��N$�'��GY��ȃ��]��k�'�Y�š̆�>�p^���A��P �����%�c0�&�cWQ��\���E��O���+��FzI���@��YL�G��E&�{��߄��Q�3ǯ0���W|�D"3��.L�ئd���`$YS5'U��)nm�%8����!5ү_]�g�=Y_ֈx�~��cD� X}?ej���'�l��(�sp�9��$ R��eS0
mf�5���m�ss���:�"h\���8�~��Kל�5��Q%���ۣ�v���{��r��զ���w��ud���u0d(*ᖻ� #���-�ii�R$H�̀a�K&6�n�,����:�E�s"����`�L&j.�����]"b�e��l��B���J�MF,[U&	��yO�{�7��:f*���/�ߺ�L��>�I\:fk��"�Uۀ+ׯ#c�b]s�J5�TU����ʲ)�?�>����9���iV!$�����A(�B���J���j��ƃHk="�����d6X�n�|r9�l믷���n��3�WP������;���r>���hʑCΗ�B tq�7g+�Q���W�D J�n	�,j\��%�Fp���Y]D�q�B��8����B핏	.�b�/����?1�K�O�f��W0�5�(�bd�Y�E-ד1F�F��n--�	3�K������cƯ��[=)vI6&�%��XF�G�'�>�嫻Ń�ৣ	|!sE���Om�.�xy�y�BY�l�D).e�INޮZ'o\OIՑ���}�EP�MA�X�p�Cg=����g�֚]���s���N#.�ܶ�ÿ��Q���?�*�	@ͨ��!C�>*�:!/N�I��d�tם\�^s3̢Яa�E|ǡ�V��M���hX�F3A����<�6����l/~��;B<֢�U�=oV���1h��_�q�NH� ^�� �D�ޡ2�$k~\���5��*v9;Ѯ ��|?}��ӊ8hrfW�Q$��3��D�G���@B�������`���Z���'m���2ePo���j���##��K6t�ə#����˚}�R5��:����;�(g���ٜ�k/�{^���`so��%���=Ue`=�)@�vt�̢[ma����2t��x�Kz���U#�D��$�W����j6�=��͑WJ]i���F��e_pI��	-У#5�Gذ�n�'4��1I�Is����E����:��_p��`��u@ѡ/�	<���V�f�bU�PQ��X��T�7��v[���sRK�����n�i�)����E��r
�3�!f�3� �3�i;�m�;pW�)����K������ ^��w2r��A�
�_�og�bُ3�)��.J����;@a%ȹEy�7�>�b/�RK��R�;J�G!f`�������[D��R����zmF����Y�ey�a�=e �����5�~����	��_����5&a�6U�x�#vlS��<'Q��)���8x���$�s��Ƥ�(5��F��!����#w�XZ�Q�Bwp虪s�=O<j��N��!k_�yq�*�!~(E&n�l<����r��W����2��5B�zmG��&�0.���v��]5P>�ٻh�T�	Db�A�V���;Z��g"�2rhBb6������^pyJ�5ΊԠ�]����9w����ɼV�[n~���8Ω��]ĳ�5��tW��Es�ؐa��k���[��)�>A �|x�7�B/� u�/�b�q�,:��\s�Qī�z�ݎc_�iz,��[�ȟ>!��.]�ڻ�F2F�Rgآ����E�Z(�8A�0}�k΀��Y%���6Z�@��8V��`�i�y����[������5�'���R��#���(fDρ2��]!����直q����iC&������~J��<�l�b����0<�H.���]	���L�l)}(���\+*�CF�%xq�k��ǞvvӽV%r�2�ͦj?}ynUY�[�����$�LoÒ����@럹\�lq9��-�M�z�\���P'Q�b3�:LJ����,ċU�� 8j�!'�R�ng7����
��^���V�b5����l���?^�ƍ���f�zY��^Z����Qp��4Xm��k���3�,|FW��Á��uhW`��W�H!�T_���tP>�����Eg8�(�O+���2�(N+���XЎ v>8�C���f�E���Y[j����dշ�.D�K�E��V�b����o��e���C�*F��ͫ�M���r�Yu�� ��嫗{9k��W#Xυ��Z��ɝkG�%�G���07Š�1�~��vUg�����t���$=&0�F��M��}��\�}o�7�#�w���Pw}+cH~�Ro*`��zg�\��ΐ4h�`�y[��d��(7O3��m6X}+[��Y���0��
}�m�|�o����`4{�Q�[Nf�zYD�xf?�4�cs(�h	8� �@	�D�kpN#��Hv�� Q,�bYI����G��$SQz(l��r��;UWlQ�+��#�H��5�(�@� ��2C�>/O�H���ApTkݪ5R�ZI�.wY��
��;�9�Ŏ��_gK ����+�	��ʾ� i��G�QIUޝ����j�1�����c�W�h����@��+�`	`�'�2��d&4b�\i���r���A�+�d8j��ݨ�Z^u��9�b8/��	�R�|*�L���oa.�5��E���P{����	x�n)ݽ�X��$�!�g.�}g��#���Yqt��.B�(Hw�� ��h��?�"Z�0q��C�E�PMb��>��/o���G���Jc�,����>�P�Y�hݷO� f�Q��Խ�Xz�W�Lm�a��Q:g�A��/�2�� MV���uTm'�$�t��h�"��>���\i��D�e�ePmi��X�`�F��Pk�z�XdD���bP[vv$�Ô����y�� �|С�Sy�x�w�D�|���NcX�Z��GF\ɉEmcK��[N���Mg(@q�������˒�ac�p�z_$�C!*C]��ē�!�K(-y�W�&��e��@�^��q��C�sZ���*�D�g!ѹ=�/�u	;xwN���z����͢*��B��$q�i��N�Fe�z.��mv��ł���Ĥ���x�)�9�_Bޏ�"���o�h� ��y�ߴ�@�v�r]�
���u^�DO6�n����5�sI��ƄR�,�9:t��=��}�����bQzj�(�;`{d�e\ǆ3��ܾ�2LԸ��?��Jp�G!_�;�r��z��k�8J�d�*���t��0�����[�x�@H%�(�,D{�t������9���x�@��H�XF�N4ѫ��mz���^�/xXx�I+ z��e��ǌi}Τ��w0� )�|#ӧ�V[���RD�o���|�cӟ̤R��m�7��(���%p�O����m���ݩ,��\E�&`#����+�ĔP�����HxL����X��mQ��y鑁��#ޣ\.B����mGϹ8� �d�;�#L���v�\%��j���>)�j\Z�A�h
rh,�2| ��©f`�y7dM�F�(��ׂ֥��w2g5�WU4��qU���H�(~��)h������\���r^.�xʣ�!���mf�ԧ^m#��Փ/F���J��y�\�:�Jr�pǬ�[?)�j ߼�����ZLN�ޥ�O*҃O�wc��g�P,ā�uR���L���M��xbB7����}~|��_4ULҙ7 32��~9S}���9gĭ:��r�`
i.{0�S�����6�ο�SW�"%��<'.�Ӱ�T@!~U��e4Y��g����"C�� ùP�� ���xf���h�L��^��gE���V� f�i�   f�������������f������f����k3�M���}�G�F�� �+P����6�|o[��&}��	�rE��>G3�J-p� �?��R��Se�<����iW��&���������X���f�4ɽ����f�!��H�j�k��h��0���s@�x�X�� d��@�%���X�@e��I}���F+aFp����S|���X����l��}y� ,����F�Rz�e�v�C� �9�:�[�(H��i�E�X���B��~�A�ϝ��@1:�T�h�ӇJC�#-H����~1�Ű�:��o����,#}:�ޕ�̻L��۞��dl�!jò羅�DE��sB����uwy�G	���i����+���dd�M�3%}�l2��؛���=�d��&�6��W!	�v�c�р�Y9��#��Ӛ�ΜU��kJ٨�Y���^�Jʌ������6o�LN[�@?S/�ϨSରh��w��_�.8�����S�����.nOGY��C���	�*�S�pa7N�	���E[Ֆ��⤍�_�c�[�9ć[�&��*"u���T¹�nT|Hq��u�=E��^K�� ��פt�a7/�f����,�I��_��@O�r�(M5���oN<M��F��yN�-d�n�D����P뼥XKV2���0ڛ�s�h�FP���[�cB<�m(�).:�_\�a��<�En]�$�� &ߒA~�f)\���f�:T��`�.I���ν)M�0~�{��Ѭ�)}��+͏W�x�@ �o����>�A������z�$P7a70���5����qL!6��e����� W�ֱ�`�*�څBW������<�����FB����֐K�Wkl?�^�W��#��ٸ�gO͍@�rK�x���7㥁�x�&���3���T�6�e�}h��`{�r�F�������gMi�p��de��?�5%��b�\v�rs1[����2$"�)Z~ �O�U>�ik
�uN���rܡ�'#�<>sί���*����Xf|+������9z�!�`R�"h_ގ��>�ͭT���CQ�Ì���3��Ǉ�����~�	��A'�n�pZ(�q�W�Y2g��1�P���SI �!5,����OA���q/�L�Δ�;,"����@ĕܢ��=���N8(���t?��������i�8Z�)��}���T>�;�9�������-��/Z�i���5���{�3��YБ��������n��b֐j`�f����;%F��ev�K��PJ�5}��ñ�l����+VW��QL3�Ֆ	�0֦�����jU	����D,i���[�����f>*K
�:](��h������"��X�]a��l�m��3��f�͗R�i���L��x��ϰ���7����7�J�zǧFF=t䏀�z�]�Z��i�y�zϡW��gp����%!&:�`��XS����ra7�u��K4�yE_�M�����VpOTR*�S��`&SV[,������-�`IT}.��Զ��?�,��+۹��M�1��͐��!u�YXV�Y�Ėzѻ(9��� �Lg��4�e�bN$���d������[c[Q��M*����ZFC���#[�(��v��l7����~��.�\<�cm#�a��R�=�B���_��<<�T$�G@��e���w�`ݸ�{�td�`k�N$�� m��7��m%��ꉤ'
o"/��NЈ)�P�3�js���:l��=J�Q&i^7
Ȕq:�앛������h���-���3�C�zt�����^�@@r�y��UR�KȮ���V�:>솰��[S �8A ��e�m� �s*}5��q�s���w�@��[�.��w�E��M���1���^$�Q��c"�;X���柪�YB��q��@C��~<蚷�Qz��GL�fm��F�tiN���$57�qV�4�_�W�Ű�nIބ;�I��[��.�� ����-��U�j,�%�����DN�Bm*z�VZ	9�MJ�S��lbb�%���Ϲ|������T4�����w�9�R�v6�	,��JH٫����6uN�;�^��[����[�\��d�� :���\��
���T����S�/�T��bm��7>�̔���Q%%�ѡc���m�M�����t�2��Dm@�ɝ��5�:�:Pe�������=����\��t�P��9�ꊢV�
.$�����k�������m�nH������G�6�0}#�GJJ0�9co$9�Y%�4>?Jz��j�_��e�a�#�x�i����an��u��]Xb7�r!�Ĳ�H5)\�<�s�:�6�1D�W�U���ok''$�{Q�֨�s׊���J��:gA�g�;�vK�XO�Ň/]�`G�$!k���%0gnP�ܢ��"��W(b�q�K�}'�yW")PN�om�����2��Y��$��j�������r]r����~i+��3y��s[.<J��h;�f%�*`�����������\=�།�+�	놨�](���}�|��#
5�(��O�p1`YvA]��8H�����+���1%`�@_��ԉ���V*ظ�PCD���K �y�K����F��d�hS��M
�� aO��y��_��r�x�5-J��j��N�o7N�[e���O�%A�h�8AƬ�"U�;7���bB����%����*�f$TV���9%��:�/btخ�QA:)H�H5��s�\��	͎��&B��63Ey�.e4ե�iP1������F2��Í��ሙDW̋?���o;�V�;�܂� z��GѷƷC��O`�g7Jլ��__}E�F\9�m�rw$K/�#��I����|F��9���� `K3�}t�f"� �6��2)^�$�HY�E0���؈=Y��[t��Z-��]��p���,��i"���B̹#�+]�r�cJ�o�i��BZ�ܹ���|بB�������,�QaU	����Q�@���&��Q�J}Yauf�������¶w�r��j�u�h�NxwX@[Z�c�7:@������g|޷"�W�!���T�\��P%¥d:o%�w��;Px�{�70׮IB�\��8rٓ�9�݌#
oI��F�V�����9EB*�Dp��S�V�$s)s��Ŷ+�(��9'2�X����	mN2���}r����	����.D�޳uKY��;�e�v�8Է�k�-U��T��| c!���ե��`����y=�u;���B�Y~
��
+HY{5,+���<}�^�g̈́F��*�ݩQ�ѽ�]�v�"�$�*��>>\�*������b��x	L@s�9��^�mu��ס�I.�[&�;ڒq9��k�T�צ�\���.��"8�o�'����_��V	uN�[b; �Y�>n��O���E%�����l��J{��Z������yQ(0{"�˛��"�×C��g�*]G/Mz�S�0�\,�4��
Ŋg����O2��6�Օ�Y��u����r^���*�i�����5����[���2�M�A�*3�����po��̌�>��!���Z�M��M1���kG0��=��� ̿7����g��0fg�9�ܴj�̈́u�s��M+v
���w�u�Ѷ;'#����Q�L��������Y{8@$��}�"B��Wl>LI��Zu1K�+,�x����_BT���Ÿ�Ζ�U�o����������� �(���k8opӊJ��!=Pw��g�둂2���)n��!�`t�b�,K��q~��J�� pXG]�/wX�g�	���B
����+���5�@���?���*�#�ܹ:�M��y'�B���+���;�(��Fj�8;j1l4�i��;y`R�W�����|4"�T�������-�&�9L�L	,��W`�)����)��8��77�"u���5��i(*\A��Y#�7{I�[��Ť(hf���OQT��E�g�/ܜP��L�0a,�a)YG_�*�R��8VK�_�(�O���@v�8��b����� }YNY]�J#6L�����dF�7��W�*g9��� O��w��XE}��zLAS֚�5�=���O%Xo� ��� vm~P�}@e�X3zeІ�VQ�n�>Ů_26]�����S�x����cצJ���j�Z[F4��eK��[��js�QY��rْ�z�l Fn1��>�mk����k%V�C���]c9�!�.�~.D����E�;`��FY���	�<���+�����1,5�a�O�)�=���K����)�����-������vhK�t�V~�#4l��O&z�ʹbB�Ҋcb��ש��<f�+�Z�0>�(������AnR?�"���I��E�Or�a�]4�gk������o��L�r/6���AN�Cε,JQ�;�3FW���žԤN^��{r���A��+<cZ�)3%�?s��O(o���k;����m���N�*2w�ф����ԿǬ�$tHD=$�ܙF����z�1�CL��O;5��� ����G�ʅ��$9�R��D����F���:B�\�b*%�ؓv[&c�$��3p�j�38�G�m��\����X����Wl�/��~�=+��۫�Q�a���~ub�N`�ph��adJL�T&(��p�	��8F#��^��;�D��v��c�V3�r��H-�X�.�~�Xz;zcL�u�����s�>i-���2�B�Q���MA�%�&@#��E;yk�0������2�s��Fn2G7oS67��7l�r��ם�O&��e���L����j�t_Ub^d��-���Ƭ.;�`/�����bi�d�ܬ�����:xά\�,_� ���Iu+�B�8Y.����b&�K�`VG^?��Y!څ�(��3�T��+F�L��w�F0qkwĲ��룀h"�'=踮r ,�Of:\.nύ2��w��~�8��y �=��&@h��Z��#�'�9txt�����'�tN��r�;8kTw*
[����1ΰTmb'��X\7��۳�:��G'�N>H6�>���t�!�>��a$/Tx��h�'�q����߮�5�-�i�^T|�1cG�+#�+���k�V+�]V����H���A�X�s�(�1�v�=��U��{~$6�����*�w���}�TMטD�6�.��Y8�ժ�-q�����o�f(����b��K�K3
�=�cˌ�a4�~Bo�D��R+����p� `�ŤI�[*a�����oS��"|� �)��@%�t��\�arN�y2l!�6�B��\�vX٪[�k�M�����]}�_��#���?r�2���mne��/�xCB0�{V霩/�Y�3,I��䉦�y��;���d�<�*�O�����"��؆����/7Y��[#$}�,rfc���n`F�	er�\��}t�M=��Ө�h�n��S�^C%��銂�q��N�D��Hխ�Kc2,m����,;5FO>82�/FN~��M��2h�Kp�\�n\���{�)f��5��%��f��?�4�ޠ���w1~�.��;��X5
ط�zVx�4�T�&t��yy\�	�nuE�g���9�T�̓&WZȏO/@�x}�O�Iw��}�����*UFad�ƶQ�夼c�A=���h��&w�K�k7��|�
}��7o���h��x���6^[����+YSA��:Ux@4���{B��U8=,a�fճ�a�X�M����.���3%s:þQk���F��b�'�ԉ��3*H�TE��HlS�����Y��܅"K�Al�#gN���~q\��,����+%�ƅJ�0z�8�fk�lQ�H^��%%P�Y��r�o�ZF+,��|�8�J���?�o�"$-:L�d9{߽��7Ԫ-�� /��"���P�܏<0ͭq��m�U���Sj�`���@�RS�9K(k��a�c�Q1�lM�S���D��X�vZ�,�8��A�a����FDim)Z��4�W���/�Bs��Rï�m��v�9ADM���ׁV����/k3�)�x�d�ۻD����� �g*c%�	�ȍ��3���
w�-D\���l�I��6�.��1��uʒ�L�9˪y������` g)/*L
 ��F��"xJ�,dг@��'�Jb�jޑFd�^�Þs���2�J$a���E���`!����E�>	�K�L#��Č�
�A�+�WMU�'���V(#�$�c�~2�=����6� �<ٌ�"�/KhR@.�fy��R&P���� �q��>*�b�u��\x)�Td XYn�
��� �a.�)+�u�'c�i-��M��^I���B��d>1E9���4�KgD���z�vE�Z��m,b~AE��=����&M9��)�)%�%揙M��Z�Λ��*�B��@R���$I$����9L��:5��C{�F���pKI�g�pM��I���c1�j%X�����Q�y~$�OO��|:{� w�J��>m�Ԍ�����)r���Qv.���{j۞TdW��26T�������K�Q�)�����viQ޾������=���h�Q/����F�� l��OE�nT���6�j�v���9g�ќ/�Y�M.���S���F��L��#�:� >����e��s�<y�<9�U)�x�@¬��7BH���y�A��!HQ����TGWC�J�B#������?+����_��@FI.�?M�B��
.U�z�N�f�����7��w��Ԉ@�
'#D�|��S=��P���~<
rAWٻ��	�H�t�8F����
��>�׹�N���/������ӯw7������_����"�G���oK�j8J1��]�p:EE�5�!IO�8�q�R�o�κG��'����܅r7�E�o�/4��=���E���b{r���Zt��ֻO��̱���`YzƎ���0{����h'����x�����X�p�T�����5��:�^4� ���)?��0�~����6�������������b:�
�q����)����$\'���������U�Һ,�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �Z-�=Q���,+�m��ư��;,�b���bQO�-�f\�f��-}-j}�f����u-�b�?�.L�D1U��cT���������{[����x���)��yS���<������� ܝ<�K��������d���q\W�	��*[�T�;�(��<��&ڮ�� �<�M��d����ª���d�?{��qq���/����� إ<��
��f����^đ�/A
���� ��<��ڮ�����{.���#y����j������q�������� �j �Z��6��哲��~��q����G��������V���}�Ц����P9d��N�����#�,S�iN��ZS�e_���ғ"9x��#��h}�ނӓ�hI����a�Ͽ���S�"z��� ��<��ڮ�������y��Q�|�􅿇�Ɣyq�����(��<��y����{����K����?QI�M��Ή����?o��s������ ԟ<�G
���O���>�Ik���Ù���П<��;���<�)�T@�#�@�$�]�������,�)�=��Y��)�����ȓ�R�i���Ж������ʔJ�� *��*|
���M���yN܁���_��D�Ej������AlM� �����Q��Q�زd������I�KR-�����h�f^�6�?CI4#[����������������������F�Z�8�����y��EE��nS�̅k�&�����N�#:��h���h���h���h��h��٧{���@MpV�i�|�=�Q�=�Q��~�h� �D�@���� ��/|����5h���y��R�|�NL�>��έO�����C�{W�Q|l��8u[VuS|T�T)���Ñ�R?i�j�����Pyg�hӓ��M���#��F��yږ����_�>���4�E����ˮD�?ZH�M�������}%LKR���Q���'�G��j�h.|j�������i��h�ŪD��������/|������-Ǫl�j�hI�������G��j�h.|&�������i��h�Ū ����yE�0k�h��g�j#[��¾�p")�M�������Eh隺�{���#[��¾�p")�M�������Eh隺�{����#[����QK@\|���#��Ez�u���KO�B"z^�]��|�s�����M����+���}U[���Y�����Rُ�|���V�~KV�x������2�KF�p���(�I�z�H�v�����C�ȅ�K��V��	��� r�*U���T�����wRُ�z��ʢ����T��Q�z'���T��%M�Y�|�X�v������%D	���K��ھT)����yp�h�j��h䋞h�=���S������Q���;�Sm]]����Kn\���ƢŤ����č������J��i����S����� k��[�h����)��ZT�R����L������ȑךPL���������S�"z��1����퇈ґ��M� ����M�|ik���uW��@��G�M���A�@�8�A-�0�|���,ɑ���/j�����t��M�����7�M�����~h���M��s�O��?�Qg��?e���{����Z���Ù#ԭ����<��q��;��N�%�X��O�����¾�pEuS�q*�޻О�]�Q9|&�c���������+�HS�bI�&�ZS�^N������ԓ��Փ���������Rܕ����q��h��j���)���,k��B�h�����,����9y���j�Z��¾�pEu�R�a*�޻Ў�]�Q9l&�c���Г,�d�������,��Вy�j�h�V�����-���SߖM� -����rQ��������6]�����R�=/��%�y�E���������������Q�P��@��*�kӑ��b��^Y�������
���4���̌V�2��[�o�֜.G�Nu3��m�.������T��ꆭŶM�(�=TR�ZYVe���&���3���g�A1Y�����Ĝ�(��]VL��w�n����q����\W�o#
?����I*�$�Bw8T�od���U��x6��W � ���ط��y|)Bo�Xv&Ǚڠ��fP{��4�1�P�a��/kE�5���<`9" ����S��V(mC��LS\�
Ǫ"�#}��6U�b����(d{DaxQ�˞�y��X�3Uy���N�]��M���{4t8����ʍW`M�C��Ø5��5D�4�#��B���q�xZ[�%ޛ���Zgb�<����؉`Wل|l*A�a�|6�(�8������Dh��NV��/���?i�3�H���߹,[<���{��WZ1j�L��$| V"+g;5bTC��P1wU⇓���@:�Z_]By(inB��h��̏\��h�
��P�I�u6�S�^�W���� �e�p+���ncϤ��c�oS.N�t	�ȇ�#�]"̧Et�k�%K�zh�$�z<%#�8���D;�-�=�<�'TP�'���S���~ u�/p��^���U��Ʊ"��}>��<w5�[�ް����}4kP��*��F �N �庖�;��'�Nu�?����I����y��$�2�e�S�W���"k�K�1K<!ִ�l�X!+�@�X�K[���JEerYu�UO$3��ܨ2 CZ	Js�a�9�
EE�-6{_d}�B���S��˚�~yk w�ּ'2�i�{�������\��A�\lb�G���Y$��*JO&2
������٫�C�%�<7D��o(��{t�b�U�?&���K��b���Q�k)��ނ�'����h�Yk�M$:���B~{B�7p9h��!�m'���{w�@��U?��K 0��@�ċ/�B)���i��\�q�"�{
T	천��E�)�$HP�qg����-6����I��o�O"������h�ft�a4۹C�\��JN��]��W�����,x�����Ɉ�-L�F��v�ɒN��m�6(ʋ�����
�IT��	�;Q�,Ά�
�w�^��<=�_?� �\^�4����Or������LT���N*�s�4?�c1�IN(<�u�U�M�㊛�q�0[yˢuh�n531�ĘsQ��{~;�g���d�Ҍc��(C��IX�Zb�|����z |W���W}�6o�SP99\�qj+���5+�r��_����J߹����[������PGKcݟ;�'��ZM��e��c	����R�]����=�����zn�/\�ꤙx�a+*�m�t�E��V:��۷'4��}�mo�n%���\�CuY�u8k��E���t����B����n���3Y;�s�#"��)��� (�JMi}�7��%k��Fi���' pn/���a�E�7e��eEP��e�M=����/i�V���-|�r��c��/���[�J�W��2�.'ݷQ6��'��<�����3��(Z�	���$�m�;7b�/`S[ۿ�y�5wa<\�,�@�M\��o�-�A�}��{��d���,��}��"��RK���T��n�J3u(��9�O���JPY�`�`�͌\	櫖�h�E�iA�j�Sm�,���	�%�\f�ݐ�o:�g���S3�j���]"���܇��m��d���@�T��\čjvب!����L��;I����D\��Gd�������4�VV�B@>�=P+���*�n�m��c����E�lP��4�цʎ���w�����j������1ec?�q.�����l���Me*���t�^����E{����f��@��݌�l�W��Yw͒���zS�W;C��1|�]����k�H�S����Y	���|��+KǗ�J��� ��.b&�}��rM��<�r��Q<R����7 }��8y�ga���n�f̾p���bb>NuAR����=��S/�2M�G~5�ZA���TP��Ҥ8�!)�Ld��Z�`�Υ��|�P�+u�r���K�18�r�\BY�?�5�I}��
|h����s�(�Մm_�WE_:M���pDڴER�%�`�1v��U����8��� ���g��>1�	�}��(���hsX5�Y����/S�wh��F~M�����LF���n���V��J2{�;�	�݄��G�KG��+��N��I�.��4h�!��_����:��K�������V4I�
�j�8�ĭB�kD�� �<'�G4�S��Ê���Vc5z�ȑog8�#r���t��O��O>G��[��r�z%)(����	[/����?X#�,���0=;ED��v��Í�w}�\u��[�-�F�PIb�\'Y�ƒ9��	��v��p�5n�w�%�5�j@W(n$�F��b�8܃��%�Io��.���J�{���W]/���=�˱��2���\j�Ԋ����"#��T9jI�����U!^̦�E����)?��rE�g.b�_�`�p������W����W�۝�1��_Q'%!�c_1j7������(�;�L)�j�@j�W���/&�в �~	G��q���H�㻝���?<=�W4Lk��e=��4��V∁^!���\U.X��O��+&����V"+�9oW���\̛\�.�asZ~��(*⎐fļ:wQ��6Xۡ=%71�++m�%T9��9���n �*� �؁���Kg|������l���R��{͈2����ߵN
�mD�^���4� 3�a.�|���j@��X ����Y��/h�P�%����-���xY�����3(#��� Pփ4T���.�>�R0���#�`�AĆ��Xo|Yq���,r�G9)���6꽘>��q��C�H�c#Օ��&�3$��7h�Ϩ5�.���d#��)��!����ڂ��fإ2�t���4% j��A�.KB�u�K�t����f�`K�`4w~��i:���
9$�g�������*z%X�����b�9
}y3e�tɩ����mE!�唢����N!ȁ}I�R<�oѳ'��F�l�W���^�G���Fab։QG��ܑ���x%Xp���W�LuZ�h�Ρ�a[;�404�5��y̓o�H<0xH���g�mOV698!Lc��-�F	QD���ڷ�>2��^K��^ܞ���-�=#��D_�����R�� QQ�_O�	!{2dQ�?��Uv$?���/��"��Ç�
�D�	y�B�:�6�DW[�4 &�×���ɆO_�}����=���-�7%9�S:rЎC�P�Wu�zR�����g�?��)�R�P][�7��AA�� ��?a`󿌕��k��S]%�Vך�ȭ�7cm���zu��@����f���=&U�hnd=?��%_��'���H�<eQ	K�z~ǵ 1͆�׼n�ET!|���ۄ8������1�詳p@���nE��Єw5��^{��%�1�Ez=}2�d�r0�	A�>��C@����TR��U�����ޑ9{���$)>P��(od� ������<;oj�θ�W�5�e���sd���n��^�\Z��F�؇�w�6�;(t�.���{#�������W�A{�Oҽ�r[��\���P2�E7ԝ�C��D��=Ԕ�4���7�̰��s������pRӕ(���!h�r�~��>1<�$ �I��3��M�=�=�=��	��TM$J���7}���b�xA��w�0F��؏�Ɏ��l���Y�a�I�N6x%|0Ġ\x��Iw���n�g��s+�snn����i=�`�v{���$�h�(w&5C�]/@�.~o���p�Lk�}Z��ѽ�p��I�z�lI�A�
0�#�d��5|����B�'�5��$6����6V��U)�mᕹ�R�)��>�S�
�����G
��R��� ��c_3�����F�!-Ŵ�~]�|���Q�d��W|�Rh�煋�Ӯ�\��B2]��*��DS��d��6�*��3���[�����A*�i���xD��S_u�l�ɒ
P;^K�<��k��D��u/��x��1��'�qt%0������'k��=�o�P�ݭ�0ƕ�7IV9��	���O�Yr�g��Y�捅e@$�a�����F����ۯN�b!���(�����B�0�e�� ?t��_([�Y>�c=)���p˖>�z�Q�7�'�.���Y�}���3�>�&2�4�\��mTg���UdJ���@�f$��1�V
���"|���\��!i
�h��v�o��%.��m���y!���v��fF���9V�*��/ۻ��@̐�ƭL���`���덻��/��_W%�͜��
'��I���k�w��@52y�e���c��Q!!��%<g��_����rh��t�ܣs�N��C�4]�:=��|��Y7� %��4EZ�� �����8�mQ��6�SbvK�1N�_�}C	2����j ��yy������)���$%{�-���B	F������*/�W�g�mI0�;�'��k����N�ƱB.���F)&OX'uV�$V,�$!t��MuĴtU�,!G��o..C��t��}�!�!�=�/�"NlИ �p[�/ס&n���0�Z	�ϻ��'8�J^W�*MR�����*DK���*2;Т~X[B��a<�	�/�a Qy�=�1�:#����Z��,F�oL��嬒`�<6֪yf�����,	E(�e�g��W��[^�H?y�#���QZ���G�,ǰ�5D�J�~C���(�s�ڐ7j�\⭤l@݃�������%@++������o�ʺj�iB{�!9�LJ�1��UC1S��zU�i���Ҧ���ų174ճ���ɵ��,�/� �QgFÃ�I�ťRX6It�)�C�;P{��HQ�*�f��E��88 V�2u��V� ӟ���#V��r
�����躞�@��\	g�NK���%)��L&�o�r�d���!b��=�,�XE��VȜE�ي���y�|�eL�O�<v��
18�]����!U�*�x�s�C/���!��p����C|D+@�N��(�I(�?���Ւݰ۶Ύ��?��:|�Z铐p�o>��q#��o�	�^��)�S��<-"U-[H
+�m����R�V�yo�Kc�	(��LQ�
Gum2��F,Vj���(�*�H������-1�8d�G~� ��dS1�`�St��{�:-s.Ah��`�aV�'�͓#����1�<_����y���((Ss��J�#�7.M��<�8����^�Y�~ �@r=��pc���=�jT�q�*}�����1�F�9���P[ﴷ��/`�W�1�k+F���D��c$�+Q�6�	�)Ԅ�N�|��>e������t��dlIbD��D�8�Z�`�+�Z�>
�c_�O�ĩ��.�e���P]�:��}������f�ޢДD�I�E�/�a:�i�+���Ng��s0����\;D�������O��L!��bY���K����#V>�v�p�s�H�䯫ſk�~��j<XOzD��N����J?J^W�f&��-��d�����Ɖ] �����>%�b���^�-cA�� ����:��H��M��<��K�Aֺ��i��-�i�p%���;�K����֋�DC�o���OWQB9	�"��z�N�>�ٱ.���4����Ϫ�@��v��@Anh+.�t!���)��g��8Bw��H�I*��׷GٖSz��^m���@��>����Re���Qad�ǒ>4��XnYneT���)1'���s��/��������_?; �2��V�"l���P��}i�����d�`hm�������ӭB
�c_��A�2��\���hSn⨺e��~��Z�]�'�f�(F��h�\x7�5=�x=�җ)��7r���Pp����
5�n7�*�u]�J6�F7p$�q�Ӫ.m�w�g�:������r�֥��M���<gpJ��?�RO��	�?�@��N�c� p����M©�a�� 5g��M�!��i�ѡ؆��W�<�1��`o;&[���\��\�O@6�$(�b��Q	GM�Y�-Nj����B/f�2��>��>Ī���coS�e�j��R:��,��������MSc�E�{�N�NZ���LX�8IZ��=�	nA��H��{Iv�Ph����t�*Ry���/� ay��|��L�۞Z����f��v�������ߑ�bP+��E-z�[��	{A����8����r��s�bO�O&��9��]@�stק0�);��8nb��F���NT���i�%�#��41�i��ݢz- 
�U�zn0S�<Y0$�:�;h��ĩRV �._sB�+�2��Yy���d�}�6(au3>sVօ��o�����6���\�<�� �'.f���&{Z��"�\V����Z}Y�P�n��1�d��0E�mÆ���}����Z�ْ��  6#_��?!@4l"�+�n)e�Kw_5'��~��;#���� �	 �LA"�XS-#�I�Q��M�x�	���B#̊|��D�&!�GX~^�ξ�|}���M0K������J��Q�I@�z�uZ�����o��AձDR�H��>�΁��A��h��D� �\�"la��h�fD�;{ZJ�C�7���r���6��01�,RO%*��؟�@*�^�HvW\�����J�{����I��C>/m.�F����n�i	��|��0(�Q7j[b��nB�<�5��p>г��M0���<$���s3��3Bn�&g(5
���u�0�m*��:-��h��%c�F/O�G�.#}l�r쫀�{�m�wVE��gҀ����sv�R�zUx!nNv���ޘ�8Շ<���U$s��Q�����~n�#���� )��5c3*�$L���0K�r�GF���N;��upEa����P^��bP#"�U��*����r}��Pb�(��W���c����}k���d��B�����&a�d?	y����׳��/|Li�7B�l�S)��&S�ۛdD/I���F�(4�]�1WQ��}����U�'�Ѥ�6 ��Q���-
%m��w_�W�,����}���%�~���"�m��](W��S�	9c��7%����1s��O?3W�R��}8�T�oC�A[�zG6��Y
/��&z5-q,���I8#����@���=[-����i;�o��%ʇ��vY��m����8 �Sg=զHT�>I��]�ZH���(�B��_�f!����>����a�@���BJ >͍͹��MoW�C��.��&T#d�5"��,��W�<����q#�]����R��������~����pd��:7����v���~@\R�G�Ǣ�j�D�7�ua%0vWa�&�3�i�ڑ��D�������y������,���j����� GskTy���"�u���}(�s��#��!b_�ɽ�n�o�(�`�������;�x�$�Pa���X��(���<u&�is�*}��c��o�B���� ��j�*ҩ^���p�8��L*� ���)��w���!��U�1f]��kl��������.�N�Q]#Z`Cݥ4P��ȟ�4�i99��s��(�KS?P�G(��uM�!��ɻ+������l����g��2f�΍�~���d�L\�b_�Ta-�e�k՜;�6���t��:M���uT��q�9�W��������P�q�0֮��X^��E�~��ǺA�(��������P�'�����GO�q\;*��y�+n�>#N��6*��� �����,�g�"�=�Mlh!O�Q;
k���Am[B
ll9sA_6�c[ ż(jw���E��e�Ns\"�)cW�E�/��G��0����y��J%��Q�67�X���9����{�R��"��}YHu8F��{h2�>)�`U�����pw
���8��G�wlSԸ�X3���G�Itd~֛� �=�}�������ؚ=s4B��)��*�;F�0WS{�������p0�!����Vw���8�(��@�/�����!����u�y'��j���y�mEN��̤@Xj�4��KX��������wi�:Ү��[ yic�Dp�ω��6�E'��} ��:��n���˘W��Aw�/�J9D�׿[G9 �Z�T�i�Fx�y'��,A��]�/��@6��:�ǃ��`���D�b
�nUB��`��2`PЏ�F�,8B������5�\3�6�"�h�X���ǂ�m9���?9�)d��̫*X�0���j�)@��w)Q���j<�ZW*��A�gae4��DE&nI
����Z�47�-�]��[d/�P�\��L4Mɣü_X�S���,�%�4P��A���]s�+�k�SX����|:!|����l��"�~����~�4�D0	����܅�o�1������bJj9�캍,g1w�;�~���|� �嚊Ҝ���L��I����k�,��r��	4�n�J�j����T��k�S'X{��� �����$���n�,�9���-K�AF�\�+W�"�y�<���?�3�-�����s������kFRq��N��'M5o��"`�-! | "���!����u6-n�@���oɚZ�r���?�	+f�_��;�pD��f5M��?�(�e_�D��:}��}dIo�Q:��ir7��D�x(���+6��DP��ˣk����v���s�o|�oPQ�\�s��)3d��J~Ppi&��B�>Q��<�����鐘�g����N�O���h 	�r�!q�t����c��{�z��mĊ}l�Wp�!8$�	���J^��5B�*������d^�5it���U�_~^��U�B�h�df+�cO4�[$�ԫؾXv�"	�g�y�y�M���5�{Tt��C ���3�g8�����V��㪃�rg����M,��b��H��wIp3�d>�h�F0�1!L��禉�b�X��zBI�%d������fvdI��A*k|�$var~�w:Ӭ;'fl)�5����8��֪H���a�R�yc�_�nu��1�����]&�	Aګr+_5�U��Hx=�x�P�cV��D���x���˔+$gO�A'i�,*l:�[1��h���Y[l혢"�J4��g���,�뉫���K⋏����t�?�R�Ri�K���,��|��%��������u�?�aD��0`���()(��!!x�J��]��2U���R��X]}q4K�tP����>���'��h��䩿@@�@U��Ky���C���Z#�O9NA߂?��\�$�D�����dQǗ��sa�#A��ήC-�:?;�E���;��P���%peMaٓ-O��	��4�WI�#p>p���Ń��������57������d��
B��H�0�UWfm$���3t��ً,�������m>��K���mю=j��F!(�����K����޳E�7i���+sb0��T�?���y���6P�#�B;�E���!�F-���C}�V��R� 6Q�6���T�7���<�E>�H)������c�MR�F�B*��G�tD����,ƍ@ j�5��ʫR�魒��@��lJ�|%ȷ��Ac�HQ��p� v�����Y�!5�ˁԎ�{@�7;|
�&р�(��`�뿐wkp��GI��/�j53�Y�HZ�<�k%]�.����3�!�P�����x��1�G�� \u0ש .�<�����4[�<�}=6BJ��p�Y��Y���z�W3J�b&� dٌ��!�q��"��iwq��j���>�j	?��p X�ŗ~�N���+�D��Z	���}C����r���_An+
f���"�����YX�xo	xR('4����g��X���v
s��Pl+�a���zo��|���@��~��)n�kL:C~�Y@����F�<�*u;�z���Lg�X�od,C-\�,�9 η��PH�Aw���BW�	���Zzr�FE��)�I^�A�"fE
�0p|�)[�q�����u]�P@,9�p!a�|	E�^VJB0?	��UB���^,{�pǌ���y��}B�vE�s[a�]�$���^�b�L����ܸ���CĂ�(�Q)����R����e`Um�w�<R�kZw�-/Y�CV7f��3�>x�����=�ւrɣ�Jc�S�=3�DHDn�����E��ʏz0_����,��5� ��	�ۋ�f/Ptsrߣ����Cժ�Ev�[99H�p�:;�3~�Z
J�8��m�J
ߙ<l���!��Z�TԺ���T4%�m�3ɯ�h�}	0I��Ff�ر���l�Mwr��#�AxIR�q�=$ݔ��u�ʊ�EW�/��o�i|�D���!?�T�v�W�Y��:��9%���(ls�:l7=ӘK��P(�İ+��W��ԅ���ۓΝ�Aϧ&20_k.$Ս���ɶ�� �(��h<Jz~g+��j7�=���A�i�c�s�nT��4B}n7��� �3��RC߉E��a͗1��os>ܱ�+VEQ��qSZ�{����o��������-F�-B�fn�9�Ū枪Mv�?���s]��gF<��FH|��m�����Uo����I�(�1-��&��%%$|�)���j�_:�T��d��E ��A�X�}�BL��q��&�ˊd+�KPh�Iv��I?63JJ�R3E.�q1�)��Ǽˬ�ס���8@��0&$B�����5DN���}^�_VB�������Ec���S�y�m�� �������LA�g��&��z����4��k��|&{���©��4d`2��֓	���L�N��C.��EV+uFOP����/�f�TT�d ����=UwĐ8{I tȒ�#�%��x9[t3�ɻ�+�EP��-O{�VnD���,�/_�Pꖬ���Hi{�A"Pm�5�h�y� .�6�1p@7@�����a7�T*ɖ{>#�7�݁F�}�ee�Z�!*�r�N�,7z�x��C�=)�gs��-������ѩB
*6-;�����s+�_mL�l�jJmu��=��5��N�	�G�W�!� nhhX/D�\(�����pf���e٥J`߁��1���U��-x����aOZ���W����K@�?oEg�8��䛦1��7;A�Sת���Yy��$ݢH��^�Q]��������p=��틠���x��Ц�Z=��$Ht��wM6%*�O��#5�Av@ �;��]Y�m�`L�F+I��1x?X>	)�%gyqu �!��*���[17lf���M�oI�����AȈ���z���d�J<Wg�����*�7���!d`����\xd�蓩$�Dz�v^�TL#T�dh1���mr�#�ʛ��I���:/��@kf��/�.L=:Rg�[&�����y5�9T���0���0;Ve:`��l,��_�Z&�t���=s�@o
&q֦�έ�G	�g��h4�yа.�~�\��#�D$nv��W��v�|�B�6�;z���B���<7�4TIXt5Q��*�� �q�� A<�9�t}䥫D)�X^z�I��R��,�����M߰W����t�Dp�u���ӵ���>����3,��Y��% �A�ۑ'��"��K��V�!Z�:���*��:��f ����9M�:9j��0R:&J�UV�J�~�ۜ����4ɢN�g\/�a��ԃ�zb�o���N�R�G*�ˆ����l ;��V=�Al?�F�ogX@\#r�&+��Xqx���
Cȯ�=�,�]U��:��z��=�+oĦ���v,�7V�"���.��sl;|7�񌳠)��ڱ.�_�g�d��t���չ�ŧݩTĚ�3j!����#U˃�*����s�h���K�*j��z%�h�`��~Ma��i�l��'}E$".R��P?㐟Q�n���D��:���3�֯O���C9�u�e0f+��a5�Y�Y��ħ��r��񸏾8�/��fS%�=g_��X��ێ"uG�~�Q��AZ�Փ6�֚Y<�k�Ȑ��$��W
w�^��n}��:ɻ#	Y�X5���	��C�)�'6ϲJ4�ʶ�Ǵ�\�[�r������n�a ��-���ٲ���\(�ox!�f�<�(���`�<�&t"��7"�~g.���H� O��]�mR\�s4)�Ǡ�j)�i1=ْ�nҗC�L(+pO�67��M!���s_�%����)Ԡ��-gV��E�'���Qmv�v�u:%�g��
���k`�51Rl��`I�e��F�VqK�����q�Y$��z�7z�I6eC�������W��!\r�4�J�J.G9z�W�u�����n�x��8�
Fb[C?��гg�ȼ���>%kM�O��c�⬩Y�&X�`�:^�������'�-��x"�-kF��7�ʡ�-�Gy�j&�C��o��4눰����F�4C��/o7O����8R���a�On���	�l��i�zg��@�~�%e�f\.�4��ֆ5V�y�� �O/�?u��)B�Z���lI�W;'*��^	+�S޷�{�2%�km?ݚA�N�T�U�Rk!t�v5'y#�I1�b�ڀ���zؔ�Q�:�cgJp�9��b#�5_��ۖ#��0�ʏ�B{�]0|�n�H�q������4HX�x�jAt<�ӥy�S�`��(#���M���z���9ې�B
\�C|<�K�UZF��6ε�J�.'�Zp��+�w�q^��&��Q`�f�
'�5����1�����'<�RX��>�_�= ���w���S b���6��]\*Y�{��<^nR��[�(�����PNG�a-�}�@K玾�Ђò[����4��}�\�s\��z#���P���T��ZE4����",���!���]�S����eB괫��z3�z)@ې�$��ީ�5V^�1*^���&?���4�vdt�N�z7���l^��(��\����l��/a�p�'F���v��H.m�D�� �Ā
�{�]~����9'S"�EEUNr�W��I��|r~(�ʮ~%� ���>��X�R��&�Y4�IAk�?:	X1�g�R�KL��D�,���\��5e�uI;\�m��_�%�����HG�Y3�lg�u�d]Il�1@��lUZM�#T�����-pQY�����Rܮ�Bxiu�h�ŸW1�@�֚����0�z��Ȝxg��i�l��1�ʃ��/��=�#:RM甁�2ݥ��p>��ߨ�w�Z��_C��ק�9�Ї�f��L:�~e�W���5H�?H�;�$�J�rӹ�A��)��.:�I�!�7��l���GGD�@�iX`A�)ov�}�	x��Lpuq&4�Z"��o�����j����|�oCK��"W??�v� ��bH�ү7ّTӛ�'UJ�x����q��r�+
�.���R���␠	X�aM�����k=�D܉=���$t>e;$l��� �ċ&�wݥ��j��ha-8Ղ�����y&u�g�O�^����뼲^���L���("I����=-���5�q�m�ֲ껂.��)�0IH^�_�0�dt�h��]a
���l������Q��f9�j�I��1�V
�%����CO�-�I�؟�+JͰ���-ߍ����,dܤ�\'Q�*6����� .�Oj���9D7��U^�	x�䩲]�#Pg��2�I��|XrC��+y&LJ爡9�N��@"��PM7�f#٧r��S��ݸ�J9:����8������K�T�w&`�%Oҍ�
�2�Ee0�'�_���3��f1�NVQ1읽Y=��3nVְ�@o��MU��gT$������|I�󀄴c�K�*�PJ, �NT���:�4�1;�(k�B�s�*9F��Cow^H�9!K�V�T�n�$`�-Bg���^�K����G��9G;�� ��P�ὛB��p	�;G�:y��e�=��z��]nz�w@T�99��l� HR*�ſ�[�(GH�I�aX�,�m�;��wIM֣�ܑ���0��'N;���ub����B]��UO�2��u6�G�Vt���~cl<`k��qY�Z�B��>a�7	^lo_m^�o�(�b5��.�a����,*������'��b���;X�xv�Ȭ�Xzh�ڽv/OG�g��#ڀO5r���Y�{tb��7��a-n%>�t`��M�A�\�y��LJBˌ��k�5Yv�1�J��p���2�>#$A (p����B��;=���/;}!S�p8q)b-u�r�f1�h�r8L��e��h�D��Z%B�N�K�ޥ�.�4�݊�Tb����1�������of�c�,��&�����di�@^w�ۮk����ˠm־�K��|D�B5[a�3 Ks�X��ǆ� h�����ע�y��?���>� �,�+!����"�U�u 1{,f����@�D�~7N�pf�U��;-r����!r�4�������Ѷ�'�7�CUcF�F��<�9�޵����{��� �����o ��9�t
��,� �g�7V	T����߆u3Ǟц���O�ԗ��ˏ6:]�4}�xۅ�����`#f8g�(�N��E�	�Z�ҨS<�le1����/F��A����C�}���!�Z	Cv�})x�I�3�p>����K�E^ �ʘm�ˉ��=�oD�������wjxx��J�B��^6I�^�㺈z��{8��օ���	�+�>��eϤa��s�B�t`P�w��&��Q98{� 	r/�C~L�Q�:2|j8<����n�&�.��+���7a�bujmi5=C��s�a)H��]%���T� �<t�,�L��u��7��en^�p|�s��F��dR'��l~�,�4_�T�ԁ��Qx#�~����M�ϐ%�����"?�<G���6�\3(����i��r{�F��h�4An0�����pBC��������9˸Qڢ)+�I�\�G��*�[�wQ��|�^�����zc�j��-q!%;�(�j�5���כ������e�M��Kt��.�3��Vm ��?}�&�}��}æ����F�xy��Q��v��(ǂ_P��O�c�U]����)��sX�o(x��2�,B�J���L�q�,���h}��K�7�Dd���� \4�#kt	cf���RȨ�%����F�Xm0	S���}�~�<��l ��U�µ�Ѱ8<Gl���&x�l�q̠��pZ$-D�����2nV��M%Og����%�~��_�
��(������6Ql��ʔ�7ČGi�;؇˛��T�Qx3�8��l�/�(��(��\$j���@����N/�]E2��{ɵ��#?�K�����1P�9aY�_ڡC筒+�ė�K�_�f&1��a3�w;7�e�6���z~���c��=���%3kV�S�)��B�h������~����{��t����;�9�
���PLF���?���g���b�ش��$�-'a�e[0�1VX�NC�ú|X�ˁ�����l@5ٰ�������pwQ�}��S���j�L�;�y*�
��P/�S� �#�G/���o�?c+�>t42`U��n̹ %@��7���dj���R�n*�4J�-]�y{ILC�P6��pJ�{���f���k^��1���h��7���� 9�6=�k��8`�vn�'p�|6~��Z�'���J���!G�T����3�����T� ~��<R^4��#�!�ȅHw��3�]�5���Y�w|��NӨeI�"Қ��r��RP�δ���NI1@+�T9���1�#��)�>r��*�Ƴ뀓OW�d����K5U|���T�#������p���!R"ZK��>�E��fA�Ƞ�3����g��C�7�.��ǅ��8$�yi\e�N�S��8��[x���g~��J�GM@�d����+.���|��@Xlf��2�e�[�"�3�Q�b�4ɥC�W�0��;�^�7�ff�o����ǼN�{(�t|'O�mB���gVH��ng�^{��$��lw��f��{K�-�G�	ywn������AA��#�}����p_̳/��,�0�B�)^�ɽ������/gX�}R��튾h�l��{J<��hŎ��{r��`F9*|˦�N^ŧ��Ig�̟Q���g��4���f���M�w�V�
�{��i,z���q�gY���;m��N�~<���d�B	qʡ��&�\�f!�����aZ�r�
�9����c��4r��dZR���r���cj ��Ag���:�Zr��{	�]�	���"+���n#� $H�2��������,�O�V�T��|]Y7L�����������r,���h��N)<�H�kL�}ns�4<A�k�w�8��'1Z'�|�}/�� ��K��}�ݯ~ɦm����U���nqG<0:2��}�����5O�W}���"�0knZd�Q��N��ƛ
e|���Foj!O�ۣưg��'��zq�j@Q�$�)��|!�aE!�Q��̓��E��P�)/�Y����j�&E�� "����z��`爅a![ O�,�Bszѩ�^`\��=ԹGWA5��
��[�q�٥k�goBͱO��0z����C�=�p��4}��ŻRلn8��b�3��ځ�np��F*�[�`D��be ��m@�]D\�!��b��}�CL�| n�cs[߹�$�����1�ڠ��~��TĪ��-��b�Lv�J8*�[[qs�ScS؉�zLE�� �,��a�p�{	<�>.ǞՂz�҇�"Ӧ��	�f\�hbM��B�/9��o�Wl�u^F�ν���=���O%u����j?4��a�8����<�����0��V�6�4���z|ذ�s�-�r����j/d��ƸZ%���Q�2Y"�ڰ@lēu��M�C=9 ?������QĪ8�C;ہ0ya�j�������m�` `�����
z{5"�T��E��Χe�S��{�Z%����N��$)<�oAU%�%J��F���?Zy���.��P��kr΁n�۱�1d?�}�z����U��lW!�K�Z�=���SpS� w<\�P��_�6�*�>z�0��/�}l���?k���l�������#+!��[�j���*�Z�>��n����&�5T���|�nmU4���w�����_����O�;81��@;$@�B��1����A3��vEw��w5V�h@�l:��b�ޕ�'l��zK����*��:�g����C:wڙ ��C�}��Od��z����[Ob��������Õ���N!$�,ټN�]�*���l\��6v���pp�M�5�5V�Y�@�5���J�n�%kqbj�8Q
|W��Z~��Ր��1A!��1!v��P}�=J����eU�Iާ"�M���H�i��~�7��\b+���fZ�����L��,�{���v��r`  y:����>�f�mM�Ø�Qԩ"�B��/H���\֨�����9��ҔI��M/�!�����c�t�T2��oʂ�	�?Ӫ~��}u	ʃ��]�S�]��!G\dĭd���@!t��e�	X�~���#��nd�UUc�Qb\x.���\PB�C�J�jnJA�
#��Y�r��fO@c�{uC�JN�'.i����_@�kD�$n!�uM� �^�@$]�׾3���Șs�Gˤ+ ���ωC� !�U�3N5�L;Y �2������ړ��r���q\��HFX��=�C�e�ʏq���}��X�XTH��C�$b(�T�z�Ao�4-���c zZW����ҝ�M4Iɏ�A��T/��L�7]p�$k]�S��MG�t`;��N,��{jJ�?��Jd��|�FKS�rA��WFR ��]F�%L�V�W��Ne�3�&�-k}iW����4T�X#7nB���m�wŴ�X�P��"Lv�T��>O���k����|k�/ܰУH��&���H4�����?�I߂l�&�QC A��
��ri��i�0`�{x�fb�6�%c(��'�[�Wu��W�}�w�L@j�J�ʛ��/����w�t�ĺ�L�	��G�Uz�& DP�]b�~sc\�E�3tK�R�S���Ź'E�UF�P�%����&PMG�y�f��M��ߟ �Σ5U��Ͳ�S<1���U-�*�R&Ї]T5����镴XLuX]�R�M�X��h� @��(�kB��J	 �����U�h���          m�  ��  Q�          ��  Q�                      kernel32.dll   CreateFileA   VirtualAlloc   VirtualFree   CloseHandle   ReadFile   WriteFile �  �  �  ,�  :�  E�      msvcrt.dll   strstr   strcpy   strlen   memcmp   ??2@YAPAXI@Z   memset x�  ��  ��  ��  ��  ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �    0��	*�H�����0��10	+ 0h
+�7�Z0X03
+�70% � �� < < < O b s o l e t e > > >0!0	+ h��A�!
�	w֊�.�`s����0��0�Ġ�{��+'��۝\0	*�H�� 0��10	UUS10	UUT10USalt Lake City10U
The USERTRUST Network1!0Uhttp://www.usertrust.com10UUTN-USERFirst-Object0080129000000Z090128235959Z0��10	USC10Unot provided10UMahe10UVictoria1!0U	103 Sham Peng Tong Plaza10U
Jient Trading inc.10UJient Trading inc.0�"0	*�H�� � 0�
� ����6,iQ]-%E�}A5��������T�{�|ʨ�#v� ����t��r5�d��FZ��V5O`!����q����x��%|�@��k{<T�,�o݀���sy�Q������$�i��(�FzVeZH(���$	 ���&p�1`k�+�^-�8�	�vS���1�q������	�c�Z�-����O�Ҝ^*��6�/����ǁ.y��6F[��F+�����c��s��>�4$]+.0�-xL��.��}=h6�i ��0�0U#0���dt�<�ݙ��[(M�<��0UD��s1i��?Ɔ��[�|�M�0U��0U�0 0U%0
+0	`�H��B0FU ?0=0;+�10+0)+https://secure.comodo.net/CPS0BU;0907�5�3�1http://crl.usertrust.com/UTN-USERFirst-Object.crl0	*�H�� � �υn�}~���i�����G�DDѵ�t*�2$���M[k��L���˭�W����v���`������B���E3+�n��o*),�5���6�=�6�8�B�Nx���(I<�Ձ�&E�����5�Z�dD����E�z����������R�IO��U���h����`V�<i�`�K(�̜i/H��5f�uRP����^)s'�ꙝ��P6����>>L�|�ƙ�t�*���`��6�� �y�0� ���9
IlX�1�D0�@0��0��10	UUS10	UUT10USalt Lake City10U
The USERTRUST Network1!0Uhttp://www.usertrust.com10UUTN-USERFirst-Object�{��+'��۝\0	+ �p0
+�710 0	*�H��	1
+�70
+�710
+�70#	*�H��	1��z��ƥ
�ȸ�N��φЬ0	*�H�� � ������zcf
��P 5tS�ؤ�]���ڑ�r�5�*1�;яe�N�;��K�Q����WP�S[z��̛�*�P?�
'W^Yg}RD� bLt75�wo���>��l�`xyt�2��-]�,���+s�}J���>� ����m��������xk�3�8r��e���&5�oYzeK����^_��i��Y7��,n�G� �����)/ye��;��K~e*1t��IѤ�M���PuŤ}�f�l_@   