MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �K�۝*���*���*��6���*���5���*��t5���*��Rich�*��c�?P            PE  L ��G        �   0   0      �?      @    @                     p     �^                               �:  (    P  x                                                                  0                                   .text   �/      0                    `.data   H
   @      @              @  �.rsrc   x   P       P              @  @�t�>           MSVBVM60.DLL                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ���j�i�j.r�j��j�I�jT�js�jB��j�۟jNb�j�f�j�h�j'T�j�K�jb�j�8�j��j,E�j�b�j�c�j2"�jd��j�D�j���j�c�jo؞j"�j&��j�$�j�I�j�i�j��j3|�jj�j	��j|g�j[N�jۜ�jf�jNc�j��j�ҫjŰ�j���jҐ�j�X�jL��j�Ǟj`��j�b�j�c�j�D�j�H�jc�j=]�j>ޝj��jSH�j6��j^G�j� �j���j5�j�G�j          h0@ �0@ p0@ .      e:@ #:@     0@ '   .1@ ^1@ m1@ �1@ �1@ �1@ �1@ �1@ �1@ �1@ Z2@ \2@ �2@ �2@ �2@ D3@ M3@ [3@ i3@ w3@ �3@ �4@ �4@ f5@ �5@ �5@ �5@ �5@ �5@ ?6@ �6@ �6@ 7@ W7@ �7@ 8@ �9@ �9@ :@                 �%X@ �%�@ �%�@ �%H@ �%8@ �%�@ �%$@ �%�@ �%L@ �%�@ �%�@ �%�@ �%x@ �%�@ �%,@ �%@ �%�@ �% @ �%�@ �%�@ �%T@ �%�@ �%�@ �%�@ �% @ �%�@ �%@ �%�@ �%<@ �%�@ �%@ �%�@ �%�@ �%P@ �%`@ �%l@ �%@ �%�@ �%\@ �%@ �%(@ �%�@ �%4@ �%�@ �%0@ �%�@ �%�@ �%�@ �%@@ �%�@ �%t@ �%h@ �%�@ �%�@ �%@ �%�@ �%@ �%D@ �%p@ �%�@ �%�@ �%d@ �%|@ �%�@ h�#@ �����      0   @       ����Q/�A�����p�               Project1            ��1  Ə����N��RF6� �J6y�zM�$]��uMn:O�3�f�� � `ӓ                                    	      Form1  Form1  B #�  lt  �      00     �     (   0   `          	                        �  �   �� �   � � ��  ��� ��� �ʦ   @   `   �   �   �   �  @   @   @@  @`  @�  @�  @�  @�  `   `   `@  ``  `�  `�  `�  `�  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  �  ��  �� @   @   @ @ @ ` @ � @ � @ � @ � @   @   @ @ @ ` @ � @ � @ � @ � @@  @@  @@@ @@` @@� @@� @@� @@� @`  @`  @`@ @`` @`� @`� @`� @`� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @� @�� @�� �   �   � @ � ` � � � � � � � � �   �   � @ � ` � � � � � � � � �@  �@  �@@ �@` �@� �@� �@� �@� �`  �`  �`@ �`` �`� �`� �`� �`� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� �� ��� ��� �   �   � @ � ` � � � � � � � � �   �   � @ � ` � � � � � � � � �@  �@  �@@ �@` �@� �@� �@� �@� �`  �`  �`@ �`` �`� �`� �`� �`� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ���   �  �   �� �   � � ��  ���                                                                      II                                              II                                              

                                              CC                                              CC                                              CC                                              

                                              

                                              II
                                             


                                             


                                             


                                         

                                         

                                       








   
                          











                          











                          

  


                        

   
                        

   
                        
     


                  I  


      



                  I  


      



                



      
               


    


              


    


           
   








     

      

       



      


      

       



      


        
      

  


           


            

  
   



            

C            

  
   



            

C               

   
                           

   



   


                         

   



   


                        


    

   


                        
     


   


                        
     


   


                      




      


   


                               



   


                               



   


                               



                                  
   



                               
   



                               



      

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  $ Form1 5<   �  H  0  F�     8*@   �'@     ��������    @(@ @@     xe             T#@ P   Ə����N��RF6�                                           b      �@ L   VB5!�*             ~             
 	          �%@  �0  ���         �   T#@ #@ l@ x   }   �   �                   stub stub  Project1    �'@     D,@ ����    (@ @@     @�             �$@    �(@     �$@    �$@     �$@    �$@  �h l �$@ @C@     4} �(@ �(@ @  4   �(@ ����        �$@ `� �(@ ����x%@     �$@ 0$@ H@ N@ T@                         p%@                                                                                                 �l$3   �#     �  �'@     �,@ �:@ @
  @@ �@  @@ * \ A D : \ GC12\ AJ,H'D  (J3C\ 'CH'/  3H13  ,'G2G\ (1F'E,  *4AJ1\ s t u b . v b p                                                                                                                                                                                                                                                                                                                                                                                                                       #@        <@@ ,@ ����    ,@@ 8l�_�L���&��
    (@             x(@ 	           0$@ ����H)@             �(@    p(@ ��  ��     #@ �����)@     $@@     �(@        ��  �     �fO�    Project1    Form1   Module1  �J6y�zM�$]��uMn:,.բ=MK���4���KƏ����N��RF6� w2է�A�nQ>]�:O�3�f�� � `ӓForm    .=����h�8 +3q�C:\Program Files\VB98\VB6.OLB   VB  �(@        	   �(@ )@ 4C@         Pg  @         #=����h�8 +3q�"=����h�8 +3q�   T)@ d)@     yO�3�f�� � `ӓ   \      . e x e        | | |      t m p      \ t m p . e x e        p a s s               VBA6.DLL    __vbaEnd    __vbaPut3   __vbaFreeStr    __vbaVarCat T)@ 8C@ __vbaFreeVarList    __vbaVarDup __vbaVarIndexLoad   __vbaFileClose  __vbaGet3   __vbaFreeVar    __vbaStrVarMove __vbaFreeObjList    __vbaFreeStrList    __vbaHresultCheckObj    __vbaNew2   __vbaStrCat __vbaStrMove    __vbaFileOpen       �                   __vbaErrorOverflow  __vbaAryDestruct    __vbaUI1I2  __vbaI2I4   __vbaGenerateBoundsError    __vbaVar2Vec    __vbaAryMove    __vbaLenBstr    __vbaOnError    __vbaAryConstruct2  __vbaStrCopy        D,@ ����    �'@ ����    ,@             ����     )@ �(@ <C@     0$@ ����            ,@     ,@ ,@ ,@             @      ����������������������������U���h�@ d�    Pd�%    ��   SVW�e��E�@ �E�ȃ��M�$�P�E��R�8C@ 3�;É]�]�]��]܉]؉]ԉ]Љ]̉]ȉ]��]��]��]���x���uh8C@ ht)@ ��@ �58C@ �M�QV��P;���}�=4@ jhd)@ VP����=4@ �E̍M�QP����RP;���}jPh�)@ VP��98C@ uh8C@ ht)@ ��@ �58C@ �E�PV��R;���}jhd)@ VP�׋EȍU�RP����QX;���}jXh�)@ VP�׋E��=0@ Ph�)@ �׋5�@ �ЍM��֋M�PQ�׋ЍM���Ph�)@ �׋ЍM���Pjj�j ��@ �UЍE�R�M�P�U�Q�E�RPj��@ �MȍU�QRj�(@ ��$j��@ P�E�P�\@ �=@ �M�Q�׋ЍM��֍M��@ �U�jRS�l@ j�`@ ��@ �U��M��E�   ǅx���   �E��)@ �E�   �ӋM�j �E�j�P�U�QR��@ ��x�����|�������j��M��P�U��H�M��P�E�PQ�P@ ��P�׋ЍM��֍U��E�R�M�PQj�@ ���U��M��E��)@ �E�   �ӍU��E�RP�<@ �M���x���Q�E�RP�E��)@ ǅx���   ��@ P�׋ЍM���Pjj�j ��@ �M���@ �=@ �M��U�Q�E�RPj�׋M��h�)@ Q�9  �ЍM��֋U܍M��E�    �֍U�jRj �@ �E܍M�PQj��@ ��j�`@ �   �U��M��E��)@ �u��ӍU��E�RP�<@ �M�j��x���Q�E�RP�E��)@ ��x�����@ P��@ �M��U�Q�E�RPj���׃�� @ �E�    �h�0@ �D�MЍU�Q�E�R�M�P�U�QRj��@ �EȍM�PQj�(@ �U��E�R�M�PQj�@ ��4Ë5�@ �M��֍M���ËEP��R�E��M�_^d�    [��]� ������������U���h�@ d�    Pd�%    �  �����SVW�e��E�@ �E�    �E�    �E�   �U�M���@ �U�M���@ jh,+@ �E�P�p@ �E�   j��D@ �E�   �M�Q�@ ��u�  �E�   �U�R�@ ��u�{  �E�	   �E�P�@ =   ��   �E�
   h   �M�Q��@ �ЍM���@ �U��� ����E�    �� ����E��E�   j h�   �M�Q��|���R��@ ��|���P��x���Q��@ ��x���R�E�P�@ �M���@ ��|���Q�U�Rj�@ ���]�E�   �E���p���ǅh���@  j h�   ��h���Q�U�R��@ �E�P��x���Q��@ ��x���R�E�P�@ �M��@ �E�   ǅH����   ǅL���   �E�    ��M��L�����  �M��U�;�H���S�E�   �E���`�����`���   sǅ���    ��h@ ������M��t@ ��`����U�f�J�E�   ��E�   �E�    �E�   �E�    �E�   �E�    �E�   ǅ@����   ǅD���   �E�    ��E��D����  �E��M�;�@�����  �E�   �U���`�����`���   sǅ���    ��h@ ������}� t[�E�f�8uR�M�Q�@ �ȋE�����E�+P��\����M���\���;Qsǅ���    ��h@ �������\����������h@ �������`����U��J�M���I  �U��B�����3ۊ��0  ���  �yI�� ���A�M��E�   �E���`�����`���   sǅ���    ��h@ �������`����U�f�J��@ �E��E�   �E܉�\�����\���   sǅ���    ��h@ ������M���`�����`���   sǅ���    ��h@ �������`����E̋�\����u�f�Nf�P�E�   �U܉�`�����`���   sǅ ���    ��h@ �� ���f�E���`����U�f�J�E�   ������E�   �E�    �E�   �E�    �E�   �E�    �E�   �E���p���ǅh���@  j h�   ��h���Q�U�R��@ �E�P��x���Q��@ ��x���R�E�P�@ �M��@ �E�   �M�Q�@ ��8���ǅ<���   �E�    ��U��<����F  �U��E�;�8����E  �E�   �M܃��!  ���  �yI�� ���A�M��E�    �U܉�`�����`���   sǅ����    ��h@ ��������`����M��A�E����  %�  �yH ���@�E��E�!   �M܉�`�����`���   sǅ����    ��h@ ��������`����E�f�P��@ �E��E�"   �M؉�\�����\���   sǅ����    ��h@ �������U܉�`�����`���   sǅ����    ��h@ ��������`����M̋�\����u�f�Vf�A�E�#   �E؉�`�����`���   sǅ����    ��h@ ������f�M���`����E�f�P�E�$   �}� tL�M�f�9uC�U��E�+B��\����M���\���;Qsǅ����    ��h@ ��������\�����������h@ �������M܉�X�����X���   sǅ����    ��h@ �������U؉�T�����T���   sǅ����    ��h@ ��������X����M̋�T����u�f�AfV��  f%� yfHf �f@�ȉ�P�����P���   sǅ����    ��h@ �������}� tL�U�f�:uC�E��M�+H��`����U���`���;Bsǅ����    ��h@ ��������`�����������h@ �������U��B������f���P����E�f3P��@ �M��Q�������
�E�%   �����E�&   �U���p���ǅh���`  j j@��h���P�M�Q��@ �U�R�@ �ЍM���@ �M��@ h�:@ �B�E�����t	�M���@ �M���@ ��|���Q�U�Rj�@ ����x���Pj �@@ ÍM���d�����d���Rj �@@ �E�Pj �@@ �M���@ �M�Qj �@@ �M���@ ËE��M�d�    _^[��]� ��@ �����������̞����:  �������� <                         <  <  &<  6<  F<  V<  h<  |<  �<  �<  �<  �<  �<  �<  �<  � ��<  =   =  2=  D=  X=  b=   �p=  �=  �=  �=  �=  �=  �=  �=  X �>  >  >  8>  � �N>  \>  n>  � ��>  �>  �>  �>  �>  �>  : ��>  �>   ?  ?  $?  6?  d  �D?  h �R?  \?  l?  v?  �?  �?      MSVBVM60.DLL    _CIcos    _adj_fptan    __vbaAryMove    __vbaFreeVar    __vbaLenBstr    __vbaStrVarMove   __vbaFreeVarList    __vbaPut3   __vbaEnd    _adj_fdiv_m64   __vbaFreeObjList    _adj_fprem1   __vbaStrCat   __vbaHresultCheckObj    _adj_fdiv_m32   __vbaAryDestruct    __vbaOnError    _adj_fdiv_m16i    _adj_fdivr_m16i   __vbaVarIndexLoad   _CIsin    __vbaChkstk   __vbaFileClose    EVENT_SINK_AddRef   __vbaGenerateBoundsError    __vbaGet3   __vbaAryConstruct2    __vbaI2I4   _adj_fpatan   EVENT_SINK_Release    __vbaUI1I2    _CIsqrt   EVENT_SINK_QueryInterface   __vbaExceptHandler    _adj_fprem    _adj_fdivr_m64    __vbaFPException    __vbaVarCat   _CIlog    __vbaErrorOverflow    __vbaFileOpen   __vbaVar2Vec    __vbaNew2   _adj_fdiv_m32i    _adj_fdivr_m32i   __vbaStrCopy    __vbaFreeStrList    _adj_fdivr_m32    _adj_fdiv_r   __vbaVarDup   _CIatan   __vbaStrMove    _allmul   _CItan    _CIexp    __vbaFreeStr                                                                      f� f��f���f��`f�����f����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��G          X  �   @  �   (  �    ��G          p  �    ��G          �  �    ��G       1u  �  �    ��G       	  �       ��G           �       ��G           �   �P  �  �      �R     �      �R  �  �              �4   V S _ V E R S I O N _ I N F O     ���                                           D     V a r F i l e I n f o     $    T r a n s l a t i o n     	�,   S t r i n g F i l e I n f o      0 4 0 9 0 4 B 0   , 
  P r o d u c t N a m e     s t u b     , 
  F i l e V e r s i o n     1 . 0 0     0 
  P r o d u c t V e r s i o n   1 . 0 0     , 
  I n t e r n a l N a m e   s t u b     <   O r i g i n a l F i l e n a m e   s t u b . e x e         00   �  1u(   0   `          	                        �  �   �� �   � � ��  ��� ��� �ʦ   @   `   �   �   �   �  @   @   @@  @`  @�  @�  @�  @�  `   `   `@  ``  `�  `�  `�  `�  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  ��  ��  ��  �   �   �@  �`  ��  �  ��  �� @   @   @ @ @ ` @ � @ � @ � @ � @   @   @ @ @ ` @ � @ � @ � @ � @@  @@  @@@ @@` @@� @@� @@� @@� @`  @`  @`@ @`` @`� @`� @`� @`� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @�� @�� @�� @�  @�  @�@ @�` @�� @� @�� @�� �   �   � @ � ` � � � � � � � � �   �   � @ � ` � � � � � � � � �@  �@  �@@ �@` �@� �@� �@� �@� �`  �`  �`@ �`` �`� �`� �`� �`� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� �� ��� ��� �   �   � @ � ` � � � � � � � � �   �   � @ � ` � � � � � � � � �@  �@  �@@ �@` �@� �@� �@� �@� �`  �`  �`@ �`` �`� �`� �`� �`� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ��  ��  ��@ ��` ��� ��� ��� ��� ���   �  �   �� �   � � ��  ���                                                                      II                                              II                                              

                                              CC                                              CC                                              CC                                              

                                              

                                              II
                                             


                                             


                                             


                                         

                                         

                                       








   
                          











                          











                          

  


                        

   
                        

   
                        
     


                  I  


      



                  I  


      



                



      
               


    


              


    


           
   








     

      

       



      


      

       



      


        
      

  


           


            

  
   



            

C            

  
   



            

C               

   
                           

   



   


                         

   



   


                        


    

   


                        
     


   


                        
     


   


                      




      


   


                               



   


                               



   


                               



                                  
   



                               
   



                               



      

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          