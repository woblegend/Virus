MZ�       ��  �       @                                   �   Q�(]0�{]0�{]0�{&,�{_0�{�,�{Y0�{�/�{V0�{�/�{Y0�{]0�{�0�{�8�{V0�{�/�{C0�{Rich]0�{                PE  L ��F        �   �               �    @                          ��                               � <                                                                                                                            �     �                 @  �.rsrc       �      �              @  �.idata      �     �              @  �Themida       ^  �              @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        jk�f=���j��5^���Z��Q5�gd��z�^�"�!�Ԣ�:�m<�&[�3E�s�4��5���.kǁ�d-53�*+y�p��k��VF0K��.jZ*�&�d*; E�=Ԑ�����W2v5{�J}���`�V@Wx�e0S�7Z4���s{q v-�wh��� Q�9t���sE�%��O�c0�4(�MX����%�s�jZ!�{���CH��^��7MJ�6���nj9�8t@!��g�nZ����BʴB����:����P��_)���c��I�}q6�>U���XL��׷`�-��&��u�=��U4 -b�CrZ�Ɠ~�'P�M�|:��\�2����m.4B7B�M�\�$e_�"�$���T� ljmb��2پ>vgo9��8|"}��T&�~��e5���k�0wKא;�G�#�7�0D?�Vu�cyHhR���Ǐ鿠���W
SM�F�)ť�JO	���y�n	*��68ط��Vw0�����V�$���{��5�'�h�������B$�e�k�ܹ�7����x��,��4f�7�a�rc���;j�X����NH;�Yj��n�ujx�2"�r ��_��NюR.bGd��wbC$'�m�g�8E.=Ӛ�i�T.���EDx��)�;Y0e�x,��$�����r8�e���A[v(�7).�o/4�����5�~���`{�����/�� 7�"��W��8�r�2Ww.D��"��=ݵl��a��f'������p��& ��n���k�U�Jzu�:ieC�S�_|��nz��~Qп�g�lW�����Z��B�D.����^J�;�I��A*	@����v��}�v^�p8�H�(���jf�HӖ��0\'�щW`%�.T۲1kJwx��.���?�C憲��؁ҫ3lؒ`H�B]_��vH�����LD�㖾;wװ�47�Ŗ23Y.����l�xo�	��_�{�y�xMy���zvx]6n�U�^�mQ�e��NLi[�d|M�h�C�'�ki{����'6��fT�1^���D*��Y.��t�-����T#���Z��ıU�4��eH�
����`��҈8R���J�S�%Z���'����%u��&F�G	'h�#-'eQ�*�T�U����yO���d���/T���m�ay_$dXt�Zw�� 
���=m@�Mt"��e�;��K����z�����_�V���gCѳ!OɳPɉn�s����������vaܾ�h���Z��2d1��M�����f*�C4Q��t� �y�}|���tJL��@*%<`]��f���R�[���ؚ��������~A������i���ܚ�{��Es;nJ-z�k5pn:�D�`n)�i��k�i�[[F\��.�[�.}��ms-Ya�&�.�X��&�z�`�n��d�#�n����~z�P�{U<{p�J�\]B6U�ݵ϶������[��?�ga0e%>~Y�H��_5J�a�Y�E}'��YvO!qR�ȣ�#�s�UQe�����͉2fiC7��� �/�q#��MtR��v��� ~w�vU����Y��K�H�K���=j.U�2�C��w ԗ;M��?ݬB=hW
N�s`7���=�W ]������I��Vf���28��B(K���#&�jw3�#0�RZ�"iyL5��`u�_�5�0���AV��V�#��4��L�ȣ�~ODL��3� @
��S��~D�C
��O��P�4E���<��̕��ﾟ�{�@+�>��YKC4�]V�V�k�ϛ���uX�e`�n�~�����w�����Y�#:1�+���m�����(���i_�HC���1��A��o����mI[k+˙W���_.0�Y�mc��.��#�B��4%��,��P�Sy&�[S�mr�߯~޸�v�P����hg@��rq�Xe�ڤ�Q��kª����W�ԽީG㹾>��}�l����`7����[���S0��F�~�^��Mӥ�S�zQ7��`{z����qi�|�¥Y��L(�~o�i��>�T��k��mZ�c��tR�Q��P��Ȭ7��r��8�4����ݴiF4�n"��e���B��#�B]a���y��e:��M�W*Y|����"=��L�V�s�4�WV�edT��$��>��lvo%Z��x�cJ'�\j��ʲ�k�v�l��(V8
jZ�W����7o'擲a�f�Wɏ~��Ù�bH�q���D�VT��$C�B'Y�b�.@`�р�b|x�GXr�0�QR&�S����B�{%�h�)}�A�Fr�h]y�Y7PF\��f �w����J&X�;T���b)��o�^�����ext{�:��q�-�t`M�9EF�e_V�M2�EV�bR��(&bV�=^��e��o.щ/R�4J�YP�'���i0	rOѫ�{�4�\�f�/A�~�`��O(겑�C�8d�� �:�#��XM��X��Ͷ5Y��#�%�5�A2�бNe�p����9t�6242�.�kU�{����b��O���޹xP�e�%��@ꅞ�p5E!�,q|ˉ0 6+/h�Tl>�8F�Lm�-f�>�,�R�J�8����+::�Wz��n��ծM���j�o�TrK��2�3ѥ�
#+Ȫ�#h@��,e��+(�Q$"v�"3����㛂�8�Q��(!��@���ͳ�6�(�z�	��.�r�bnu�qnC��5cQ,P������(R׿��S�:�7R8��	�dI�����{� 4AtW�矢�����������t=m�)�Ʀ"O`pa3��)�����Պ�0�Cl�͔덦���gV��|�]�}S2�^�T�A�p�[�����+���R1����O׫�/79��%�S1��QI�P��g�~�v��a(�l��5�r��^"A@�&�?��>&/v�����&���"��'z�N�(��lgJ��sW(�>��y�kkT�3��=�Y�H�w�4W>^��<8N��?��x��&>^n�{��9��-uy��O�m�B�V��[ֵ�'C����-��u�U$ȅ�2�
�	+ٽ�5�f��V(ǹJ ,1�T�M��ɕ�g"|f�V���d�:9�R�h_��'i�>�r�G��5��.Vz�a���t�Ho;�h��]k��|Bw���T�V�@��%�_zg�s�Cn��.�y�Ưu8fb�QAe�IT#	�-�����d�W>���0���!�Ӭ���"�i���*�U�p}#��8�����&͑���0&�Z������4��k��qm$]RR_�L���C��[��uS�耶8n�&��}�'Q)�}�"�a����kp?e���?�j�E� MAK�]x
�9��Y"�2�e��ӑ>���`��$�88��� ��yo��e���������kl�ra�XU�0�����7V@���	"5X��*�l�Q�?M����+�p3��|0>FbW����4�J�D�8�Bi�x��١�0"T�'�y�<W� E�p�F��N�ҚK�WZ3�u�ca{�V��4��=l	Z�◣�!����#�I��Iջ��v8�="HoAƧ��W�����O�WFG��������݌�HM%�E��_�jl{;$^A,8�Ǚیb�/�
�p%���-��T2fzUc�Ä�>��ϟ@��+���:�fP�@��U�pm����m1[��4k��3(�����k����9��AX��\�_%W�OZ@4x��f4�U��?G�KڰD�S����9��Xz�3��f�h8����Oك�.s��k3����Y1]i�z`�T׃�c]�갆}���e�W���m�q`�J�j��Qf��\��=`U�;�1�@d�ڣ\^�!7�Zʀ�y�w�}�8e�틿ĩ�:�T!�-rM�TB�-DU��=�p�H.�ʠ�2 XSUf"p&�N���m~ �"��P\j��j��3G�d��lZ�3����'� ��e�3�ǉa�2�e#�[S��ηc�8�n�Ez}}P3&���7�Cf����"������j���/R�*9��ʏ�"Hz=�_����
�O����|���ld
�Z�b8241|hr��M��vIRjB���xG[ꆑ�e��v�TT��j�ϔ�k?#�;�=2g8�A��3�*�t�@@�0	(O��Sp�%Ʊ�n_�Rf�l�]FQe�6�'�E��iK]*��]{r�n{���w�n�r��eF�l�I�/J�����ڊ���"����}8���&������|��ȬJ�Mg�7~.(�?�-Z�����Px���5��c����d��j��_o�U��mVj� ��.�``2��ƫ�ᎌ�HW��1�Q_�b�4KdJø���nl5���F+�q�p���YaJ��c��ա���(sef�vw��޿RK&F�):�%�#IH�-E��,�X�,֐��`�˙�Q�qD2<�����/O݈��O�%��� ����R���5�4j,U��7�#�f5j����א:��V��6X#J9䗊� (`����^}ԝx�K�q��	���	HX!���q�CD��E2�����V��!0B�p���Sr��s%���L����������#she*K��}7�/��hXئ�p�x�A}�/VȪ�I� 9
n��9m�+x?\[��yr
�x_�Q�W[D���S��BKא�{K�*��dX��4���7i+%#9�V��mV?>*"Ä�7��P����$z���&Z�!��TX�+�N'�Zr@�D>Y�z�?:g>ç���R�A�E�x �'u.�X�U��	]�e�N*�"t�wF�{c�.���X�L�&����QT&PWޛ	�!+�R�p^�b����Lw׌�L���'C���MQ#�߅Ri2Ie��N�-�ѯ%Q�U�Ү$&Й��y�H���P���{��>(�-�i:�Pހ%�kp��'�X.K�+;���Ϫ{T�l���`de}�ѽn�c��9��p�p����C�+�skH83U(�	��&�$�>k^Ӛwm��)�7\a����k�,h�T��R�ަB�=�@�i�h�y6j��u2u5�h��]��0t=-zh��5w�<t\`-��,Jvz[��J�n��4�П��ao}nx��0B�ݓ��>Jo�Гd�Db�v_
J��^��a�����$�_cUo2i�t�w3�&���6�90+Q�kUt�A}g������e�&6C��uJ!�&Tq�M7ɇ����8�f&��X��Q]j���7?�-��eD�"M�./u��I��2u�9����-R�)G�����)1^��$a��1�;���E�
K���2Q�V�3�}��$�x�PS�^qc����Y��IҺh$��B+�LiMK���wO��upkl��>�C���e��T�S�:�y&ԡ��G�esZ­R�υ����{�mҰ�'�Şڗar{�J<��[���/C�=*�i�xC��d>N�%sг
�ҳ��d���r���h����;�-r�t�4ζ1����8*E�t��V��l�0z�7���-�����1I���n�p�n@�o��,�H�*��@�E���d����\`Մ�� GԄ%���� e�U��[�p���z,")l%8����.DeC5����m�w��X�{���ת�����r��i����_��cU�a��:_�}�G:��~���/��} ��hm]�� ;��x{����*isPY�Q5gAA.<�K�Ij�.L���46[��r%M��ws���5��vM"��?Q�0~4 j���'���ĝ�kqqg����f�����tN���͡�U���58�]Ƕ���ᷚhF=�yR�*�Ak\�p�f(0 �
]�aZ�\mh�G����)�h ��C�.=�ݫe8�| �,��o�].؉.C�i%ލ~�9��b[ND���Xɬ�G�"�ap�29�.��/�5�<�Ѣ�3|����I��I�9�Ws#~�hLG�*��oh��an�b��y�,�� g09�9 �#Vp
��[�l��./�OA!4R�=�M�ŝՃ�	?E���j5p�]hl�>dȡ�[��3��I�Rc�N��u�5|R5�X;�{�~����x텿dCW�e���gP&�%g�e���2�B��?�phK4�B��=1)�vLn�� Kǩ��g�,�p��v�C�a���b�,��P&/�ѹ���lJ�ln��u�P�'�S��j�Q���Y�Z���cz�	�+���(p��'���0y�(	)Zg�+�e����:�Jv�d��"����R?��/�[#��?Y�	.�0�6`ɣ?�2g�'Ld���ջ�s;R��P��p� ��MP�SN?XUG��M5_d"������moN�M�q`�����)̓�n��0t��EhPV_�F�[a0b���B������e,��T{�:&�~> #@ �djE2�ț�Y�3�3y繽��$`���bںW!�"�nWX(�_՗��BPo݊:�|V�7Y�Y�5��"0_a<$C�����)���%~
��@���H��P�,�H���L��U��������z�^�&�{qZ����0�%�-�(��Y��sŉ�t�R2��� �==!�	�K����3�_�S�e{�h�*�\���X0���~�?��o�ݎg$�
,H$�����Ӗ�sۄW����Lb���'�彵������!�B ����s��q�l�֭4�Ԫ��; �Sr�۪�G.���'�q�J�>-�$�nj�kL�������tn(=�2��A��!��5��ݠ]zW�)w�U�m+W�l����)��K�];o*��1s/"�N�p�
��^�?�^�SDZ�iKݏ?�KwKEҷ�	cx`Z�i�U�ŗ�={)"��"1�t*'����t�B�]T��Ʒ.�A��mV�SҺ�{�^�c��@�� Q���}��B������a0�k�u�r�ְ�5�:�z���0^YQ���q{�@��M�W�&�i62�I���/������Zb����r��@:R��Is��ms�߸m4,�_n��dh8s4�I�(e��*�+��o&�H�&�;y����H��%��%��b���d?�\|���a�9�Uo,@�~�a���k�i��=܌k`���p5!fM��n�ГL-qw�O�eh�ZU��-`�+�����J��n��A�����5>d��E�Mw�g�Q�{�U�&���Q.���3.��a�i�Z�z�ti��C�3Z�X��5f��IY�^&�{ޠ����Mdj_�ee&�T�U��}yPᦝ�86Fb�I:`:�^j�r��0؂�f?j�-�G^j��uI��_W.C�$�=
Ȍ�f1C0Ɨ��$]1�OP�8�	�G��*�A�MD'ma����-p���w�9})���m~%.@�8Ng7���lut�|�V�Yf!�=8'wtz�;T.[�Д���.��d� 7��P�:�����+7s�~Jx���"d�F �s%�y�P�� ��[`
,�ȹ�O���:��v�(��xa�-�<��糩���8�!�\���Ԧ�R�7��ﶌ�0��hR1g�V����A���DV*��V
S�����|b�ɗ�2W�,;Suh���W��
6o�^�s�m����ҽ?��@8��N7N�YI]�_��yn�'g��y�Ԩ)�+�a�j�yIz��G�0���%��u�oP0#x6��5�~ה��^�cx?���fU
��<!*mz�v��z����Ё�"���G��c:�b��]@ǲ�ǯOg�a������c	��K��pqX�d�ƫR*-}�'@#*'���5�3g�Rf���սWPR.=�/�ݾ4;"�o���-%/wf>Ǻ��/�é����c��/Uu~(S����gh@C�B{��� D%8���9߄��m
C�]dT����,�V&����5� >�a���(|+t�	�Ļ T=`/c҇�#4�Q[�x�K�/`ݿt5F����U����:���\��9a�3�4�T?�S�D�(�6����a�^����S/���D)���T����86��+��&n�L�_}
M�%>
J���]>9f�������q��
Y���D�4����H߲x7Bw`b�F��c���Ny:S��D�Gf3��R_&��T��ޥ����e��E��mJ\�O��Y**��Ig�R&��Ù�OmW1e�G�('G32�R�!�`*<�'FQ12�n��qJ�����Qn�(���f-<���#ߥS��j��C%�e��؟��j��S����%�8R!Xg�Qlo�+G��׺����k���F_���!��CQ���p�{�[{.~�4��bao�&��!�xd�L��~p��Zsk2�ԅ�kE#TH��f�R�W��E(mm��ɳ��kS��Pm&I��U��W�.V�r�Ov�Ya���Uڥ��E��25k��U3��O�ʦ(](h�fۣ�6>Xѕ�r�lf�Sa�n֛} ��O��d���<3r�k2ң0��?a�ȴ�DJ2kR~�j鮐j���o��h8Th�~�g鮪g'�XQn�(Z=��ǫ�JW�����NH-f�Yw���Aҽ�Z�:�E&���l�濁b�Jz�7إk��y8LIz-�\9X��2�-@�?M��Z���\�-a�n�~���W5��5^�-:~(�y��;Q�&�Jrsڋ�]"�Ad~3�_��x+�)sC�^g��q@wD(�e��֧���@0ةҒ�/=���J��m,v�o.]���EpcV�~�g2���VY3��j��bE(�E��!_(��}p���D�;T~:�n)C�k3'��ôP-b���w0��AT&�6L�QF �Dbn��� ��TpA(n��=&��W�.Zk��?��4�e^&/�X?�Q�n�������V��hFR���nO�J�z0�H�:dE)�H��&��M��H_0�iR�+C��0��Rxr��d�1�������W������p�}AFWjP�7������w�^��wnT]�^�Ӑd�Y����r�W?��4w��Ms���PW~�9�1��X�RZ�SyRFঘ�z- �p�Mz���ئF��]������K�����¯��OY�QI���A��m=��QU�[���hc(�C�^�T���b
�Ĺ�kәzZ��]�W#%z����tPdD��΍7��*C�錼9<���D�Mx��fim&�r�%q�B�y{98P���' qQ>�d�4������X�Wu~O����	1`����Q�w�c�SH����/���(�1�HP9�ֽ�����cDP�kR^Y@�$�j��
��R&9���%J+ņ	�l3�&�i���l��{�4���,R�ѭ��h�V������[ ��o&sN ��~��J�e�����K񕦇�Z�ml^f��� c4Ї�s��Q�9Gx��Oݼ߱�0M��:��m=QQ����١g�&mL�pAB��-�tŠ�Yc�R�M~^J�ZXMx>eXI�@� �а�_l5D�XK��0���"P�<wZ�#ݔH�& �e��F�o�֬1|�H�v��R^��*�]�z*-yTC��#�.�f�զ�~�^�wwk�.XhA��]��b�]�k@���-�����x�f̈́��^<f��:���J#��Z*����<*	��"��.T[-�|8���|eW�>ok/e�\n+D������4��[� �p5̑A�.L�9x4�R�S��dt8]&-b�۹-zO6XMc[��R?)HM���cn�Ï+�{tߙ���Z�r���U����Y	��c�9@u�~b�,�>�IҮ{jT0�/���#O拣���kP]��e����;�(��4��X&z�;$�抄�m��z#_(�cٱ��f�O�V�7�(7w�L>���������*g���`�P��Ed�C~eYq�"�Bs���h/�v&�o{Nʈu���`Y�[hXM����SEb�+�VO�^\$+8=�ۍ6R�_��a�s����km�4 �U����Uo�nׯ�4�4� 7�����r�K	��?�nC�R\�H��2+y5��fM�*�[K0'�A'��F�g&�X�&���#6G��N*쪎ҭyj�.���)�B�(`�@��y��3�s&��?o1Κ����7PZ��R��"�P�R��R�C�}�JJ�c��Ux !嘝ٮ�_�xyo�ub���k�yN�Rg�8� ��`�C@:�N^AL�/OnZ1�a����!�,�<�"4�T8`z�X1Gº0-v�%.��v�_[��Y�t�ZS�U�ff6��x�b�3�|Y�Cc������*f������!� ��R`�-*t�7{�[�.~d.�ѩ�׆�� FFeC�Ho������\챠Ya�i}=>����p=��:�8Z�0���)W�S�j���pCe����0�tIQJV�o���o-��,4J�~���DB�&@l�E|�4My��l"5]�ݑ���e��Io��fa�����IN����v.Q���:7S�ޯ�3گ�ִV���"1h��?�͚=t=X��@��A�p�U��'W��R:��+o��AØ(�lB.B7cF��t��7O	^�i';2�YW�jH�(/.<C|MHp�p?Ү_jOIA���Ex�����_�g��k�E�w+m���f��GȍӣdY�)���!�	{m*(����d�,�":>�E�$�?�fx+>�<�V#E����"�x�����J�Ƚ?^e
'y�v���.��<w�<��Z�Wf�%��r)RY�cĲ�����A��ڻ��5d:	�*���"�Py&rA60e��˯}[��e�6�e�6�f%�RD��
��gF��vt�v{�,8�&&���D���&�Q��Vd&��
�h~v:������v��z7-�U>M�r�.U�-�tO�G���,Z@���&-w���7��^�e��G�& *i1���o����A���[��w�CR�<�%�W?p�a��e�h6�,Bn�+�#X8�J��V�W�U��V���]��Om�p;�~n|�u�{�KH�j�I5A�Xu�`��c,����ԕ���]���쒬&*�y1���]�#g���cP)�f�>.쭁$w����M�=�h+*�^�AuR&Dv~���~��"P�k�e,EN"�!�'��H�SPW} �΁@S����^���*����D��$'�aZJ5�7f�I@����1���*��A������BF�D��mo^�${i�k��^��x
c%�~��s�^f��ߨ��_����Q�z�]�XAN:�5R�B'�8UF�;Q�͘�@��U�GS WR�焁��=%�A�Ox&B����b�a8{%
H��uDWB�c�����w
�`v�0��w����зѩ��T�E�G����F�laN���(�ڴ�lD%�1l�z�t*�����N�e	N�!�E�.�<�1�wR���8%�)#���eY�$�5)z:��1]v�3[(౸0��\��G��Bԯ��	���0�wH&�m ��~_}E�q�.�E��\	k(�>c��ޚ�/�O�=H��.-�J�{�o��3t0��S'^�l��웑�(�dj.Y52p�bs*)sƻ'�M��h&a�:1i5?e��e�8�"uۘ����wAB?���L�[��q���(�|y�q�;�B޻���O�/��ۿ�Ń2%ޚ2�~;���H���;�k�W� �$A^N��;硅�w�CH�Ц�iV{(%��,}�.@k�uk�QH�:gN�Gj�A�,z�w�J�߇7�I��ɵ�'d�v{�Qv�4�2�1�V�.���xet�wtٕO7�U���(X�1��L�l�=2W����ңBO�H���S�dO+��^�'����s�Ǥ�_�����(\ ���n&$w�wK1R�O������*K�
��<�Aɍ�@�^�]�-�=9�H<i���(O�ȍ5
okwR������RnY4�auc�Ko٘�h@]�0�Ci)sR���
2h�S�Pb]W#m0����V0�]���č�1l��%ƕ0��?�F��/����`8�E�w�<`Z4U�_o��:�X�m����I�>�?���/~��V���o��Y%VH��1�-mw�^(�p���T}X&�(��^��b��|��^|fw"ŏ1ҙz��!�3�����2,»�M ό�'T�4�!�o��&_%q�n@>��ET�T��͇�ډ��CzOj%�ԣ�c��àF't筧?�&ꅿ�h�\��3���s
����W-x�2w�[X�F@�p�}�ɀ��S�� /y�(<���?�!��0�,:�B mǼ��j���U���]-�l��m8���q��ȂQm2�� ��r����E~gQɍ��$���������Վ��Q��i$��ǚ�sG)�3���'�7k�>%M+;G�NE[H3�omS�%����rw;��G���L�V=��.`R����R�M:J92D�� �.��u����a]�g�_~Qz4�����O�D�c��9�O8�>�n��|
�?�笰%������y��v!���kW�5*3*���j[z,�7PŌ�
�Ae��2_��v�X�J����B��lF:�ux�C��8(��~�P�v���;����"��y"�����Q�?W4vu&.BxM��y��\��pT�M,.���:)vKA�+2^NO��}ds�SZ �b>�X]���`x����. �0f��DYԌ�ބr,I�S/k��Z�&����HXDr��z&���"��.-g&z~�݇��۲q�3l��^�&�X���������o��7�}qj.fȱ���yA��Z�2qI(Lw�����M
��9�a�i��|����G&i2�����u��2=:���ֻf�L)Y�*U�ɹȑ*�'P�a*�ޕ�I���1!(�d��yqJ 6�=7X�uU��(�w-8�A8�7dn�q+P��e8�Rdj�q'T��I8�-df�q��F8�)db�q,���8�3d^�q3���4��AZ�O�խ9V�bB��O)Ց>VlB���U d�tq
>��Q82d��qD��V81d�jq�J��Za��--P�t�8C,��w�`��@����l�y����C"��y��9u@5uJ#		�`���8����³�p�D45{J�@�z�[�7��9;@�X	�������rquR*�LL��!}j�i�`��mU%���:�̝���o�|R��7Q3���ا��/Q	�f���󥔇�$/?kָr�p��&l?h�ʧ�@���cR]I�S�F��&5o.<챟�A>��Z�5��ϧ�^��l���&p�	�<`���A3ľ�U�37�WK��n;��YI�;��n����G3�Þ���w"D��wVD$~e1��O'�V;?6��*�Pz�/;,�?���~���|�cA���w�k'�B�&ውH��R�2�*(|���XݑHPP��U�:`<����N{��� ���2;߯P~%ҷ��wQ�{^T�����rwi�gZ)UDyK\-��q�W��z.G����y���|�QhmJ��l��{N�I�jA�a�.��R�}��	R���!P^���L62E�U�D{QC�"e#�D��dZѲ����2V��-�w�=D��э0�;;��H/�׹�d��2��If�u�B �Z��0�O	β���L���.8@dU�q�#�3x	-(=�e�٨UQ��2FA-Mӝ�"0o��aO��ڟ��J�ƛ�0��<k�Qt�Z#}ei�0%j�"XI,5G��"���Z롗���[:�����7���۩�m�S�YNiS�
�Q|�}�[���H�SW-�|Z��`�j�����X@���y��)�S��f-!�>�x�rc���@�f�y�:����-&��!Ҩ��EQ��wp«а�%B�U�"뒡��f��8ڄ�Mb�h5�p�\���X��*7��7^��^Y�YE
y�Mz.qR.Ͳ�����6PS��92�醤��*�g;�+ۦ�����U�:�H�j:a��_��&S�й<'$��Ԍ.6�Ꙏ#�ۖ�R�^tb�+�����Zu	�+X9��m�B�J�8j�oA8�
��U��c��(��Z���'��,���%���$���h�ۍ׬P�Y�*V�z�_�/-@_b�xG�)l}כS�}]�G�m)�D��J5O.L�g�KN�����H�05vz��~�ojj��(m�̶Ca�d_��0\5ۓ�O�k&{��zb$�`��BN��勮J�7Y.ZAe�xފ_T��v,�bV1��/���ckVD5r��c'�5o	O2<�+EP�Q�X&�R[Tw��o�PQ;���o�#:�p(��'
;��f��U�M��Mr����.pC���_�����i*�5_5�-nw�0V��Э�N���^�fT��Rǎ}��9)%�s5�����si��l?�k)�Ѣi|������qЛ<��g�/?q���?�p��<xд�ıS�N'%"���uvM_%3;��)���4�񩊩n_+��������S^l�N�ޚ5z/�]�5Rj�w�rʁD\��n�{
J�'�Y�1~���E9^J:屍wǮ�R�c���M^G�����(�g�뿪�B�t�x���K{�E�X�`lx�Yp�4O^f���l01j���ᮈ�dCu`���ڣ��N����ґ/H�g���{v�eG�S�-5x���j(�S��|L�5Pv�8���[�[���1T��{[����}VG�l�P�Σ�Vc���>�3]��Z<�E���qߊT֤]��o�b��{;@q3nM6�ֿN�צK���]ϻo�)�ݚ�g���apZ-�W`�i~�cOr4�!�s��)�3�`*�(�D���ZЀ^��C�$S�
�QXB����hUЫ��wX�!k��.���x{R\j�Q�$���6�NL%䄹�>`o+���w�:��f��˞��|�ANU�$x��k�&Ȫ���j�m�x'@z�2�3�B8,R&كAnXR03��aI[�R�H�섚 ��6���/Ro1I4��2�.��,7G^��J,c��Rr'n��e-��/0m�����"�H���i�<���ya&�����*��aD��t?�.e��뻜c��y(��u\;�u{��1��'���H�Ҽo������F�e�!
��P���l��'M{��&�	>�V�Z��,�:Pt5nc�d"�"�e�(�A'}o��T���BD��VYF�l��ָFD:+O�Eq��T8�Ε&�c�R�b	�|U��̦a�#W�4�V��f������w_(�X����/_��
��:'!Y�A��S*Z�+�;<B��(�"��=]��g������g;�Sr&|b��ڲ}쟟V�.�"�YM�T���Ho�I݅|�A����QgW�O���
O��_|��I.����U5+@}sw��q�>�҇^E��/UZ����;�l���aO�up�C�{�Od�i5�"��`��/C��3j'CV�p�r�|��ֹF��;T��\��Ԇ�V�Y!�?��ǉ���+*!w��#9���#�lL,l�o�9��H�t^�Z�m�k�E2S��KC�Ԩ6K�fd"6���Qd0���cN��3�I[��"K%�->����Nr��>��WpnoZ���F�N)�f�GW��d���V���l#,i[npvklOI�%�L��%c��mE7����Ҵ���eh����ڼq�4䯛�4����ֱ`�I���K�k�S^�^Df/ާ�~'�K�sU�!nB/�����մ]����G��S�|��t�X��,S��5�g�|س�eM�~AO��V�w3��}&)aJX����/�T�	2"�w��m`�n])Js� 1?���uӓ�R�IxZm"iq"�X�zm�Qr�,�	�R�����Z؇�)�k��o�vB+,ݫ('�^�~��ZZ�OD����p5�y^%�Ad?��iEX@o⩤�(�a��v�$����G5�D1�]���[c��x���g�?��|[�e�d�$�`�.�;N�XC,$%*�ܗ��s�uT�P���[pi���D^	��h`��}x�p��Q���l�f���?^�%��Ef�C6.Eޫ뢖@Le��>�wd��V���7��I��&�q=��Z�zZF����Ev��� �x��;g�CDx9�@,�[I��(�?w��{̅GU�=��q';QD�}pL�q�E���%��Y=8A�`�AM�y�0=4R%p��ǡ�gJ�.�G�eK���AcU�`U��1ՎtO(�ĥ/��x:�J�JuK�`�.�5�͆kL�� c���셯����N�uF&�}.�"f��p���/��e ��H���N]%�$iӫ�H�M�4�PJ�š*x?DB��?�HO��F)���#�$��A�j�"s9b�#��/19s��'�0���]�oD���Z�����z���i�9W��yǔ�*n�,�QdW��0�����b%O����J�\U<��=3 /ŗ�cP1�voXe�c�u�N�9-�ݙ�I��X,ɤS�v��+@21�-R ��h$xA���nfGV�w��vw%��5-��5z�F.Fy�������MԤ1Iuq�1��̿�1C��7Xr���Ih��[�wL)% *��/3FZ|F�֣�����r�A�܇E�g��P}���Y*gKAUE�U)�HW�$z��;� /~�#D:��)�_a;\R���S&����w�0R�|�&���V��^��H�(�X�J��E��#1��"kfe2�X8����M���Nj�|[����ɐ.}"�(��|C�-���F���S[.mVN�gGgU�߹f�0��!�^��Մ�@��1.[�y>1���;�~�|�vw�&]�%β�����[�Y�fZ�����R&\X:�v@���X�O�P�Z�h�+�yS�9g0!��:�Ҧk�f���؇2��Z2g�1Q��9��:�UN�j�)yO4��_fYD+-�B��bJ0��(�=pA���y�1��lJ�Z����Y�����a�nW4e�)Л㜑Q�^�I�^�W-�}n���Hy@�)��fN�'���R�&���x	YS�a�]�rCxny�WW�'E%���eK��:x�M�����rǛ�i�f�1�f\F����2��w���R�&e���yC4Z&V*�2�U��1)9�IX��^g|�E�{.��2�M�=O��[r)L�%������V��.��Tu�C&�_�U�i���w�&R�6����	`U��$�>���~[��,[�a�N.�4���R�}RA�KU2HTgҗ/[ʝ[��aPV�y�}"Ɠ�*�����_�S9����?�ぐ7��K���+�Wy�����rfYz*�r��W�^��MS��8��@�����Kr�PB�%�+K�3�E��e�;6V1�)-�}����[ir*�2�U��%ҙ'12\B�U���mR�&u��r�A��v?f�Y}�N���n��hz)��h���]��X�S��?���)��2��w��i�fVYj�fѷj���!ֿ�~���RA��A�y|N�\bޞZ"�v�N5�Q�V�x�U��Uy�_o�Hiz*��B�[`'q�7�u�Y&Sx�q͝�e�N@�*e�e��;��:"{�R�[�n8�`��x��wR���Q��[R���Q�w�V�QB�uD*�Z]�[�>8�b�2թ!�h>�~f3���۫-�`~T�7�.a��B�����O�2�h�)!W�.�G�)	U��WL��5NU��S"���Y�)���H�*X%ac�)�cŢ��.���>w�y�_��WR3��A?�\2%���*��A��l���"eE���{�I`�r\o�Ĥ{^N��n:YU<�C��@��=�[�_ұ[��iC'�m@y|^�Ƌ=.q�[�}
�v#�)���b��ʬ�s���%/6�W����|sE�-��s��#�ZA�/-�}�Ϳ�R)����`"}�CZ��uY�U1��ӝ ��{��;-��|E��[*'�O1ݾr�ٷ=�蛲��_ҵqg�R&��XZ�.g�%���V�ǧ�)�"�<v�y��_YoV����;2ֲIS����Q)*�1�RZ�UM��-lw�l~�n�F�i|�z-4~"�S)QA>*���!��C�M�tЇ	�QSR�=���Q�Y�RrRD��lD){/Cn&��ƚ7s�u�Sr�bYz�w��P�7W�6���/�!A�׍0ũ�bU�%�P�f�Yv,U���'����,��=��˨-��h�+�&�ヿxB~n�_���l9s
c/>2�x��{eO� �e�A�R�?�C�XgD@�}�2���=�/��c#�^��wj���<�Vl\
��S4C�"^f�����0����.�xC��<EEkQ�_��Ԛ7 ��:.*x�1_<hHX�{�)D�#�_$T	�
}�Qˉ��F-d�{JN!�4�-On�0����ZQ��B� �`A�F�\%.�-�`
ؾ�G_�B�C��<�R&����J(Y�o���׺�6��Z�I�8����R�So4X��펦�=�2<a&sHtR��CR�G;����ٸ烄��ťs<\<QF�"zl�Fi"�IJ�z>�A$}������5��9|�lZ6��>� գK�d[.�uц?g`�k��8�o��覙9����`GD<\�7�pŻ�Ć��5w-hj��Z` �	�Ct��U�"���T����D��{.��ܩ�.�l�ET'c2E!$뻨XSOO�%������x4(/��|��3
K��D����e�|EKz�?T��׾P	�*刵:xƔy?l�#x������WB���_0��	����H#�4=�矗$B�/�����N�_�._�bQA�S�Ӎ�d��z��2=��3
�-5�<��k$��(еʷ���ױ"��E&	^۩-�����M^�d\n�F��=�=rl�߽�u缱|���8�JcZ߆)�vh��U`��6����`R�w(�ǵǯ�n�N�y Q�*C)6�W�zV�3�W5h9��c��;����x�/�x��9ȵ��/5�}e9w-9s4)0�wrw)c���~�]L���n��i�V��x��E>Ÿ�B�����9��,أ��g�9H��O� �w�T�N|~�X�_woYd���֡������U"�V���GA���_.W�u\���3�G���.~�sh�9K=X�$�bUd���̬Pj��Yv��[��?29�̘'�]aZ��d͓_���.}��q��?ٮ�f]�K��a�&"-�3���Kə�ded������A�i��]�e;.���V>W^g����{��`d���c�PU�o"��+�z�T�~�ӊ�mM2�R2��^��Cz��B�յ��zZbwѩ�\h`��GM�N�7����D�uX���[ºU>�9@nT÷�uٗk��1�g�9�#ԦԼ�MK9�D�5�v*���~n�o&�l] -�}
��kK*.�ť��髉.屏���B�l�P���*���W1^�b�C,�2�#��S7K��Lr�ƶ��f�ǥ%o��Q�>R�#Y�1[����c:�tJ
ZT�x��@��B�+s���H`g�7j��)��`JEhk9�#�ʎK�,��-�%E���=L��*�!7"�V_���T���I�3�Gwa�!�������c�G����3�A�yOR\����U��0X��%R�`�����ҏ��l �x��hAM���e̊�\�K�ϼ����º�Y+C\`�P ��8G�i@.=�t��x�^�Fj���������Qޜz5i�"��>������	0)������\����}ct=DYR$��mX�\�1�o"��J���h�j�% ����R~�*�Y�s�$kAc��8=�$D�p�.�8+r��""�����āvRˌ�(����1?�SٹY��Ȓ�4���� �B�y�e�>Dj�v��(����A�
��ܑ��3��lGZǶ�FK���-T+K��=d�S�1G�=h��ۛ��J$ʹ�L���S�:��Gگ��ך�ύ�	�����s�� �.,_61�<g8:�mW���Syz�����'hX]�� O�^��K����3SV�@J ���� ��)�%Uz
N�t ��JOO��|mDwh3���L���	r���7_�}w߶�pn-�NZ��V�;q]{xw$ �V#���0D���},e���u��F�%�w�F!����Zi�y���.@�������m��(�2:���, ��h�`1-���#c�GFq�����ʲ��_����jS���B��F�kn�/pR��\o�'o8]}#��p ��E6"XZ@��y8��4:��G��]��u�3er���EZ�(�Ps�?��k�W򫱤:&��S�q��c��v�N �\�E��X�m�PB~0�I�3���K*�`<J�/��uD��I�����=U�}b(a3��!H���>�dKD�
��Oz^�$.�D�Z��P���J$�(+A���w���zZöQ��c쩢)c&�|5F��?F�Hb�SJ�!�	c��%��=�o���V�r���&V����a.jA���:�j4��4��#	��Cs���E*'6L�8��7
��^��#i��Ԓ�tk�._Y��ێdo���sR�M+7�.��7V���;V�e�Lx?Z#	�"Su��p�VMd��#�Jup� @���ޫ�ފ#�P^���� '~�H�7q{�7FA�qQ�ZU
؁Kp��	�?
:�+&<��A2|J�J���]����J�<݀�.9��ј[�'�:x��O%���傞_�]����z-�A�f/�$��JJ���噜^��
[Y�u���(���΃<�S�H�j8h����l//(�����so�V4͎3M.�}@˞uf0�"<��"vX[hB��Ѵ}_�H�R�g��
��@O�����s�M=��-����+�1)z{��1m�1.��[�w�9cY%V{r휓ό�����VS��q������u�
�� o�{�z�֘&�~TRS��CJ����0���Wk���1��Z�Zy.0]S�W�!Ɗ�~��11�
�lG�8�Bt%�{��xX���'BPX(8�r�-� U���p�饗~Zq�ힰ>@�/��&S��D�Z����@*�<-_%�{��<����NV��>�cV�L�	�*5?�>�ć_��RZ��7��t%�QɈ�ORR�x���<چ��_��k��?x��b>/Z�^���x�{v�e/vB�e�E�վ�%���c� ��;���%�)�~�8|�o����S��P�ڞ63Qt�-A;h|���M��ژ>+�"P#�bB��H1�z�_�:����n��G��=���m�m(O��8��dn0�Մ���zySya����$l�b�ڪn�h��1���y�(�9�Ŵg�(�IJ�BQ���F�Tu%��j�d����q���
��рc�^�l�h�w�0�S������ܑ��{����Uc���T�'?��}���i�ֺ������P	Ԯ�]����{9d*�	}��k��4@����2�U��J�7=�D����Ҧ�&_*�-��ĝ��Η��w�RrJ���)z�|m�rg1��Pᢒ���F5Ҳ��T���9���!+/��.|RwȪ���%��._��kRm:�.�ӈ�c�1��NĄ�<j�y�ʣ�b �S�Tr&yp��d�±�Ԡ��O�P�t�_�b�+ks� ��d��Ay_D���!��^�0N ��1�T�eeL��^��E�:�Zn�Q���F'Wm ��<�x�/�[���h�z�����j�O#	^��P�ա�;7�m����y���ԓ#m�g��.���� =��([�.l:)�4�Sp$��,2��4�T�0D㰐{��毚�/�0�/QK�bc$��,�^|;k�'�B\��b�h�����"�1?�zq�V��la4�c�6�2ٙ	U�O8gf�b�4����k��ެ%>�R�C�.𩥩�p9��.��	8R�j��U�n�.6&�z}R�
�E��Blm-�.(�J�'�w ��)�yl�9x���Y��h(�6n�{���k����	�sBO>X�)C	e�X�:IJ5eVK�:4�P�p�ȱD�K�:D�`_V��a�f2$_�l/>��P -��ٙ^��$�c&��/e�냕'E��{.*��	g^�T(��������o�����U�	����QB��ò��u�2N�L�C2}b���MZj���y��_ǧ	�qhKfz��-����lB�(j�W7j�x'z_~w���$4�_6�:g��=��$'�t�޼�=s:-�1GB(�JM�q�P2_%�	��p��vv]� ߞ(T�Jd�M���0b$�l�OO� T.�=Xs���Tq�a� �f�Fo���me� m�{yxqsd��� ���ŕ�"p��;xBk�MT�u�=^)T��z�N�>-��Zjg�E�{I��˓�(��}0��(�?tQc�Bo,�� �xa�AZ�De2C�HQkj��OWe��?��=�V3��v��F���H&df0�=��?���A��1r�9&utC��X��T�"�*Ԯ���Ƞy�/kU�OD����FOD��z.��Us�V���	��߰Cc?8LD99���PYU.�t@8(Vs,���/فU$7s
���e�"�.{��hw.2;቟/�%�*^!��k��>ޠ��՗l�t�0�z�x�KWc��d
�D���7¨O�L��45h�}������I)�{f]�C��H�.�tD�c������МP��h����A���Q������UL̖�9�0dKױw�$>�,6���[2�"�0qE�{hW\&hӡ�/%�5��ʦ�/�9~���e�����m`���_��{s� ��2PqXYs�UÈR"�.b���i�9��w�(�/r�=�n�U.n�X*�B&~ng���ڦ*�w�eS6�%E���Gi� �4��t*�IR)1�7z��t1��!��!ô2Y��� �o�;�x�7���4��#�:��Q��cG�";���
�<�$rK[���Ж�_��U�Q��b��x2�)�PƯ� �(2�Zc��S.և�{���w~��%������vQ��C�˗��Y�?�i�  k;lj�6l��"U
�ע��gx�*`?��LQY�ս8bU�!G��%P��wҵկ�*��
���%++p�
x�����u�T���R�u҈zb�SM?��(2Qz���NxJ�I���"8��7))G���c���Лw�n���z��緟��MM�{�����q$=fS�_5s7TQ+:a���ⶱ��4M+�2�D��E�m�b�&@qb�x�i�u���o)%��k�r�e�{���M�#�q�Ɗ���"�(�!Z��˩e��V�X�O8����+�zҸlp����~`��&�"��R�2�����FF�7�_N�n1��a������c:���U8Dn�rA��P�q�g�\GXKͬx\���T'p�s�Ѫ#�r��&Z��=�Zu%?��N���.Ж��3T�>��<9��r9�/��Io��QX����;&�
B�Qq�@�"Y��'��5-���v9��䉂z�j'�+nR2�nN�[�e#�.᳊Q��j9��b�����:�PS��:]��\����!�"W��s�9iZ�1�E(	��,�����;�>Q�:��0E��PҒ��#'V��_V������Q"�����>g�3�A�n��]���E� ��):T1�z&��gb
"��|��ay�]膣�u�g��}�'D)�D쩷�R�1"T|xN�[*߯"dzk��]��Q�P����S��m8��T��9��"Z$�V,j��܍۱�KC�S����}@Y�i|������k!�Pe�X���x�k�UI��;7�;	�<��~J����|_ª��~���0�C�2�fA�&T2����Я������Mr5m��n�g����.�ӂu9���2A� b�q��/S�	.�=l_=W�ĩ�H��@�T�仆��d�2&�|5j�{`@������������|%3�o�;��;�,�q2|����=�cA�M��j�jJvP�c�Kh"U�w'��n[�𻸔2決�,��T�0zDJ�/��:c�6t+���n�T�u����B��{�T��GK�����٫"h"r]�B7"�����ۉx�s���&�-(� x�r���Կu���.mB��Af��&�~3��z�Zy����U}^�!�7`FwL6e`�n|X��p����D�#?̠$I$�*	c�P1ĥ��-L���s\[�3�k2m�}.m�ݭ�{�ץ�N%�Y�yg�ͯkT
��=��[���-���}�c��/�'*?a4�����oQ��qJr�iY�.Lf�.@f�93�X13VX%$f0)����睚��C�2a�(�k�m���Qa�*=�+A�)餯Rr���zǟ=�ǣR^���α���gy�Q%8K�y��.���Nb�Y8���7ې]�h�4q����G��8�I~�10�����ICD�#��|��JNp��+��"���!�5�t)(�'�szECQN$�e�#��y�A=x� �e���*���0�������|\Z�A�R���%2�U��9S-ԭ�G������c�߯_O�_E����$G�}zi{JE;;BR�j8�t�|+�M�Q�B��b%��>n��
.��X�)��n�,�)�8IVc��p`!%+q�T�Y���z��/�N��2����5�B�q�o�OxJ�4�A��&�[a�&e���a.E��Ze% *�V��?tn&����X��)�z{!��w�C����9���qД#|=tX ��72�WLR�����:@��b/ST;+5o$I�E|N�~eښl�d��H�<��hg〞MA�1f�����4�����-Y;ʭ�O9���70D��·��K�'� �Ҽ��w��1뇐�V��������,[R�u9J�~E��V5.��p-�� H�t�q��R%1���Iƥ��XKw���VT�=oU�d:M�~�luc���on$2=
�h�?r׆�Z�m�ZL%��ǞT^��怑+��Lt�T���[��V�fۻ�0mdAB\8�0�Y&��ɮX�����(�Zʥ�Œ�q�ۙ�����e�	1�B=q�%Hi1�1d.}���W�G�̲��H���d/�����S;%����Ȳ~�%cQ���DUh��@�cAu"�.��
�<���*"H >��X�,��66!#`�_��3RWp��zF`QV��g��9�=軉1k.n�S0��d�{C�)=�{+��-'�^�b�9J.���n0�*�vS����5l?qo :�w`��3@���S��!���2S��V)�#��"C��%F�y��?*x�C��IŦ�9�T϶����Į@��Da,S�����O��?���&����8>UfzOηV|N�b	r�>짺���~$�� jJ%b�z�	�j;SD~;�W�^�jrDx���z����FR%�!��ݵ��/�{�JrkV��Ӓ��`n^�J��;`Xx��ȝ��R?io��/���9~��x)�7����X�I%��R��1�X����S�Й�N�{�b4,5��ޗ�b��B��(^O4�A,z{���J��++(d����:;7��*I#�`�R�[�I!��m��.񉑊[����a�e���������+�I5P4�ζ�"���0��W��$��w����?Z��Fa58w\��#��ba[�z�������r?xq���.Լh�;�{�w���Jj�~�����rhki�H�c�s��^ӚvkW!��m(\U��jS�&[!h7ӗ}���Ց �L��_����#`^��]$���HrQJK�����̲�!a�$c��ҡ�Xt�Q�$��s��X+KU/�fd�[�����x�_xT.wJ����x/��Qv�,=��ݽ�a��j��Np0�jL�d�7u��3�l�Ai�>�s�U�l��I-,�qP>���75��C�z������^D-L�5����@/`���tE�p��%F>�	�ɀR��\���m���z�S��r|O�)��f�F�	�8�o���,9�m9 ��>0%x*�axhj^�E�>�НG'�39����h��=�`�|v�=���}�5N�Z���o_�/�a�@=W0��k��I"�`�x��$DlI(�GF �p���J�oD�*ۻ_���w�� ��n�*�H�*����}l8U�����{d`�"yk�\tħ�=�����O3U!�n?r�u�+������f�+����(�,h̭'1ᩬ�[���	���~r�\���mP���@%���6�AR>j�V��A��F�;��}1t,�62*��m��h���M}��h`��SO8�z$��cn$!@F��J�ݸ���ort�[���=H���7���J�}�u��5PT|�& �2s�&3>5G�/�ձ�9�T̩%�s"6 +��^���Y����[��u4us��2q�·�{��N��_Ѝ�J�khF-���8ig�wǻ,���s��(l����p��p#��O�qDN�����%"�`=1��a�.��c;eJ@8�'�e���יv�yn┸�s,����faV3c�B���e%SM�4�&��z�&�|$����&`D*|w*o1d�/�Յ�Gk�yM�k>"Da�8C���8>N�n<G�
��6�ug3z~՞r�Z.U#7���~��,q<���f�~*�D��Ak�.F~�*VG�M�_��l?����u�l�	/��t
��y���"���q�Э��4Ω��DEkN�!�3���'t�RGxð�<�����q�י;{b�4=�m2�KV��b������҈�g�S+��\b~�N��E�
�;�����-
=�Ī����-.r��e 
%�|�QIV��ܕY��. eh���M�@A揘�$Y�&���y��QN�e��QEhG���x� �l�$��$����w2!5�9��S�﵃��_�a]�:�&$Ǘ�uj+w��ڱi�:l^s�_�.>�Muw�?��n�SH[�kƋ{M :�� �Q2�i��w�1q�`)�������kp	����zb�D;�Ǐ�?��d	|�m������D��y>~v\ؐ�o�r�a��3�;��,�]�40�/l��u&Λn�C�omBN�Hn�J��������/�)1��1G���C�="h���s���%����q�P��s�&��}��h�8�`f+�|��wX�}�M�ES����}# ��nf�˲��g��FN����.9�_�{l-�_7y��kI�`%ɉ�l.� G�w�3�]q�)j"��I����mH��m�	�-}m�U}��xS10.��t�1rX*��<GI�iJ�F�|!�S��#pq#TV��pS�Ď@GvƠ����	a�%��]8�7��@^����-�mL�oܙ"�t6�c��m��U��:h�M1�t��S�+��A�q���Db�3�~�LN���m�������KV2N�������\Y�2��bedY^&��xP^��Ϋj~�'�h�k;&�s��>R����=\�wr"��ex0F����pw�Ur��L�.��yBQ/V����R5H̑1o�>ȇ���������]c���ۉ}w�Q�������n��x���PEm8�����
�v�'�� dX�wq���h5�w�V�K����w�-��)�SZ1'���6��Vs4��>���1z��@Hv�q��s`//'���q�	�i?��F��WG�@�f<��'2 kBw_�e+���3��e�ff3<f�ksK%�i c��.6�V�2��i4��|w�|���ZrB��kd��!�m��|7��e:��>��g"����ݵ)���o���	�k�u6Lq�~W|F�o5B�E1>�Z�K�"�6���.�J��aD�xTd���c�ɫ%Wdb��f�,�ef���=�,T8��j3_��[�?��7Y�c!��p��c@"�r�4&0*0���]�����ءr�Jp�ށ�:�������}��x^R��Z恲%i��3�.Dt=�\z��v8����O���R4�������R�3��32����<݈:�^������>�C�8�����*�2�5�Б*�/u�'�3kN �5^��N�46|i_���*B��6>n�-~��2{*o��u�m3��f|�v��>'��o�6+p�S����WY�����R�R	�x`���b1qq�ŷj�&s1��wЏ>3�*���^�C������><s8h�U�"3�	��L�'f���a���m��-�;L]�G�I~q|&���W������dcr����9�q��J\������-�~ �aA~w_�������g4�kxɴj����ƣ";d@�kK*(�'���|/�#~���K_1�r�um�j�2�O2��bϹ]^ִ�kv�3�V�,�8/�Um���yZR$md�tj�Z
��<��ys3�ՠ��o>���n�a��mJ+��Oc|V��h`�_�&�;��K鰽Rԏo�˓��Xdg1�B�I�?xT�	{j��O^4r4��X��A�97ӻ3F�W��_�.X:ng3��Չ�:aL�eO��}M)�3V>�m�P`*���XWY���O��3���X�ߝ���yCYc^ ��K�p��&ј�@���s>zk8Y�Q��2j0}hfcV,��٧u>&NM[�l�BH��U�5�	���Y��c��s�~-��?��q�6�P7��g�o��/ l�c���	��A�Vha�,>�{�*grj](@N����X�>h����/:Z�M�w�ں��.8�=R�@0��k.�i0�q�~�򈸘�y���BI/�Kj�q�t��Y��oc3>l���en��Q�-y�w���bcp��ٵO��T.s�9��

��> t~�^��ӥ���
�,����U��V0k�!\�?��{o��K��hg޾bb~�r�����\dꁤjP�F�]�%Cε'��9�j sH;�e�I�?M.��Sr�g��CF��?dR�\Y�����Q�M6�>4�ebg�az�|·U�J��tN��"'V�X�]sƊ�R��u��$=V2��R���1�s&M��p���pfw]o�u�7|�r�\l�h�3خ���=�:�Ӣ�x��a�MF��$�^P���2����/��Q�>k2��'�kRd�w�F��y$Z*^k�/k&�(�u�_iV�`db�����*7�7GD?�22Xa^�����O�b��d�N�&~5�dO�p�p�d�5�k7�p��:s�����7��bzVs�۶��7��b{�r�
�Ǣ�s`)�m�	1�!�	pnR	+���������CH�+�~����xk�y�!e�E�h���"�#�d��2v;V���I~ٵ�(J�* ��t�2+ɹ�O�����a�{�q�o�o
�g�G���7x�*-�g��m����#�k�c(�0+���q�n։{i�2�6��|�.��~eoܕnCq�"�a�}g��3Mn��vX�ѣ���6�e����`��,�_"�Ww�d�Uɋ�n������eI%�'���1����#�|������N�5V�vKbc&��,�^n?eY&�A9OF��o��|[�����z�"�a�3]�-CO��Y"D�f&���b%eB���3|�2�̩���9瀧ܷi��	\qo���22����(~�����*�S���6�@"3�nc^e�`h�_�C�N�WvWtx��y��#��m2��e�qU<x'�m9xb��-�Ypc���pztv�%h"���3�a�&��4���M��)F��vq>���V|$�e����BE�>�3�At<Y��۶w��A�:6E�jy{���&�Q�����s�p�}�� ��>\L.�K:�x���C�KM�1��TL��A��oP�xl:w)�nX��[1J�@�G��<�LW����h6���"�ٶ��x>6r,{^�t�C�Og�`�ùJd/,�/�R���5�,6Q�7V(��5��L5����_s��YHʸ�Ԧ�HhV{��4|g�=�I(��	C�D�~PN�X�����L$5������E�h^�Y��;�Vao�9RP�[w���q�����
�t�Q[�F�k}a�����:)81 XV<�[4Z�/�wp�B�b�/+&C����X�5���Gr󶯱5g�+4^�R��o�m���Ub�jl1u�5�5~�P���K3��p�����ѱ��rI}8c}a'�*,��ΰ���C*�����h�l��n6�u	��I�Z����HPL�)��A|�F�-�{Զ;�r�e.�Lf~פ(�G��?��׬���d5��c������*fE��,5Nu,/3~����{H�]���C���J*HxCF�/ONe���#k���Y�OC�ՒGֱ"��}Ä�(��J�PJ(s���������t��3U�8�ɧ}��4��7��mR�"dPf<~�(0hd]��i&�g�Wmol��󿆜*P��Mvސ��VN�`�6d{�G �/�[S���{��[�
��↡^W=��8�{2��%���$<JCP�tx���j�5���I)2�fcX:]>�#�-����WN�3���WR�(TV��$�����	����7�π���3�w=j��x�@+z�VX~x:X��f0�Vی�i�+��ƀ+�A(e)�O>�ώ=��Lh#o#�\�ʓ�QCr�Zz�Ti�(��5_b�@c��S�"���5�[�����I���X�P��A=r>{J��ʉdPڦ�#HDZd���`�MI��.�Q5U�lb �qJM�?��<l����׵~���g��.Ѩ;�/<��2X`�����1r:�Tr?<�M�#���I��`�fJ���eR4�Wq�b�/%FaE����}�7�~�vT4q�{�em4�qb؛�����ҼVP����Uj��5ဨ5�h�LZhD
<Rͮ�f�����8�����%��φ:#:ޏ5U�&#�%�I8m�y��-�TAe�U`r�n�ӏ��8��7��X-F`�Ũb��04��K_�g;T�h�px"cћ�%��wqz5%B�
e�����E��{p�ؾ�R�t�S�i�U��A���^�����h�W�J�0lz�hJ&��Ih.:Y�B������pCÈ��� JW������H� S��j�~���»ۭ���Ӝ)5z&�O{԰���Tݣ�J4����M��Ϟ�l�q!/%�4�tnK~'.	VT���q�n�I^�3�ȔK���+��'����R�Nk���G&�A�G���.'��$�H:��ORA��'�ղ�8�­�2ƃ]�Oy�б������9�Zi��9��܂G�xuWd����7թ�U�{��g�A�y=�|z�?I���Nh>T��;��:�� ��Jt]��pnʓ�Špnm'g�Ā�/TL��Hq�^+�%.mVda^x�B]+~�Y��n3��(<���I{�Sf���{C�T��j�@>P�L���w}�u_-L�l6Oi:�B��yS}	���g^{ˋ�1|���Z�}�/X�؉N�2�G4�sI%�\�(9#�m���m���˔&0g�>.J�*h4���YF�G�=�;x:+����ѥ�g�/� ��iR�.�kb1e>��SH��c�f�m��{%���h��iS���`Z�g j�tǃ�Oũ3�9զ7F��e��N.7=��-6]��!TV{��FҰ��;�)rpB�.]�-x��ۻ2.s#�%�V���Cj����A]�j����h��>n��D��qx���TԮ����~���z"׉�B����l�6kx>L��r�`�ː1 �5`&3=)/OB~Sft�9����"`3#z9z�����(:#f;m����%�5�xM8���R�v!�^�EC��%�b?)���o�v�s�e���&�煃}��X5H�z��y�/�V�G�9���&�\���ä༗+�'�>�&�W15���6I�c��ltX����#��Cf�x��Tm��� �2�,#�B%xR�q=l�hi�����O��/��dzM���O~E�`�`D�1�w����2 �Ej�=�8XB��T�c�� �*m�s�#_Uy�f�'ԉ�'��;�G����c\�wW�&`6%+�$�Α�W�|��x�K�]$����~nLI���v�#u��7Nrg��XP3JY�lij4���c��]PUթ�=?�@R{�q�.i�	|=��M��'��	�t���M.qctEi6��yW�Ur�[��p1�����x�"�z���^���_����#1f��a���v��V`�X`�J�1�*��*XL� j=�=�佤崗<��(9�_[�*!�2(���
hû��Qu�Å�_�d�	+L#������b�f3����v����9rб�H��ت�;�B��Ovd�V�y8uk�AJ��5���n�P��BUf��o��A��7��t]�5�Q������w\�����2�w��s"��Mm�C���q����H]�Yd4h���bW�:�1��hDg*xi��9��'�&�M����+�$���O���^?o�!�HB=����H� �5#q1o�C��Q9�q}S�NU���
���G�����բd��`�^�l�:Տ� �lS{J�u&����KԤP����[!h͚�d�r��I�;JSB%���!Qi�3�}��>ꈅ�� U┐�I�2L�cf�ن�w_�H,1$:��E��ҏjZ�iO��Ԑ?�ewn&֚/~�8����r75ՕP�"e��Ļ����m�$�M0\>����^6U�b�ς+�)BV��t��T�m����?[1��!8���9Y}<R��D*Q��93`�<1�+{���1T�V<E���B�& ���N?D��ӻȨe��Hk�&�dGV�a�JV{E��~��e�U�A��t�u����e�>9�k�\rǇ&~�x}�),�I�S���0���W,�!�7$R�;���i��Т�௉��
�,�1)�A�FK'ˣA�A2U	肟�=)��~k��@rt��_:���{��#{fCp���X��Kd�y��7��ΥNT�e�57�K{��`G��QD�7&�P�y�z�
v�q5hJ>���B�ܯq��m��/
�{щ���>�?jE�E:�ǨR��RFH T�y����L���蹼�]:�n@�'�'�U��%�P��Ce�g�J�YP�X�ާ$�bra�b&�4,��H^4ę��Mه>I�Eײ�����(iV:f�U��TCĵ���Z�_~h �C"�^�������OHM�Ihv�-�uW9e�;��8+R5~����������,���̊b�k4��n>L�=��&�|�S�\�x؛%nH>+�JZ1�-G3xsH�0F�?B�_k�A[E$��.]RpzZI,���7��j�Y�r̹!�VA�G���~�}��$��m���J���ş��%iV��59��gw��y���}�'��v��TK}�}r�nY�"P�^Ell��O��. k60�=��i��%���sx�o�u��;�-�k��Rb��(:i���8��b)��o�$��g��a�ΜB�)��5���{���^��MR��5[~��?���6�m����m��[��sp�o�D[��H�5�'p�n��`o\!�����h��w�W%�$������,��(���<|Tu@��'��nv��o� 4���5&�bh~�6JCe�����5~���`+.1Z3,�9��w	g?c-iG�w`�$r�,%�>�"b 9�o���qJX�a"�5wr"8@�� �����a@Q��g��7R�����8U�aۍ�:��6,%2&����Q����ٱ�n�g����!���/�<��� <�.[r�Em, ������z��^j�VN>T�u���y5C�e��q�=�t&x�1	ߥ$}��#��FH��r ��IޝMi2��j3�*e"��D���3$z�+��g�ѩi7֡#:kr�*�ʪ�>6�Z�7�&QeL�X�P&1^S�s�3#��KN��[���W
�ڰ:�Ζ9����Sw\˛]=qVC��c���]x����-(�TVH�sD�.{��X���4�
r�7�͈�Vx��p ���1 u�(]��f\�5*oR�p��O��&O������q(���&D�	�>q�^HC|Y�A�?��ev�^�]�!P\�~���_�bbग़u��A��C��y�8��6��ˮ@�9��-2�վQY=,N�D)R�s���׌ �����O�.�~Ԩ�
1�����ܒf����j>���ģ[ts�K�?o�a�w���������ey��pS���2�dp����X���Q{�r�T�t���~�A�k�!dE�ԾO	�e�T̪de�	c�
��/	��x@`�� ��F	�u�C�����:�
A�~?^��V��bL�_�\�A�_x��j3�dyO��Oɐ^_�P�������ญP���`]�QǮQ�t���Y���O�3?���r�d=��g�w2f�s��݇_����ͭ�Uf.��-�Q��E��֧�=�m�Ҷ�����(]�i�e7���G>FmW�V�g�&������e���ꖧ�=fm��v�ǝ�M��(T��4��. T���&HDJ,$(�K�&tzn;���XB�/d̨0PЎ凓{H�ႏ~���f8<6~3�v�4�x&W�\�p�X
�)A,�.������]��l��k��j��i��h��g��f��e��t��s��r��q��p��o��n��m��|��{��z��y��x�vD�"n��̯V�lM��
�|�_T�x".�R�V����i\�����}�J(���'��C�a�I�fN?ce-
>0Xq��^k1Ύ�:Y�Tsb��E���26_���h�+�7�Tr����$nE��Xn��v����� ����
��N�m�^O�ej��^r�\<:�y�"�!�Py�[#~'����<ۍr��lMd�I���>[A|6�LF����چ��Ǭ[y
Xʹ�Aה�5�x�S��y�.��8sʗ�A��T�%)�s��椃������Y�ř��6
��fS�υ,��H ��1z=%���;
����YN�g����j2M���d)���i>kF��TzA��-����d�=��2��k/B��G��9"w�y���QNq�i�}�}UVq�O�D�"�V�	#��M��k~G3r�r�S��X�re�˷�
��	;3;��B�G����G�~�UOӑF`���;��iV*��Sm�k4�^�؅������	U�����#L�qF� ��N�2�~�1-�1��b#�%���_æ,�>�Dɛ�T��������A^a��'!���t�>@/�:jny��[�z4����c�_&U��7�J�
7{P��s2�)\�䠒Ώ���	z��:� _����I��|�2$������5����#
6�::�M����Å�&��|�bF
j7��z"&�/Iz��X�y<�����~D%�7~�!�b��iۊM�?\Cd����D��]�8c4:a�4r��ҷDHq�}����J�]9u�.hP���?u�KVQ~��.+�VOc����.y{�p��N5
��F                                                                                                                                                                                                                                                                                ]� k�     ��                 P�  �             y� �                     KERNEL32.dll   CreateFileA   ExitProcess COMCTL32.dll   InitCommonControls                                                                                                                                                                                                                                                                                                                                                                      !��Օ � rQ     �    `�th�    XS   �8�ua�E�-7 G ��������=@�    X% ���3�f�Zf��4f9u�P<л�D  ��g9t-   �ڋ��^ ǹj ��
�^L �jG PQ�   �    X-&   ��  � ���Ha�  l�Y��h�ځvArv ���?�v;��c1�L&����x�^/�E"��d���u�T��k5�;Wa�+M�.R�%���<�2CclJP��u���v;��c1�L&�X��`�t$$�|$(����F�G�   �u�F�s��u�F�sO3��u�F���   �u�F���u�F���u�F���u�F��tW+��_�G�   뛸   �u�F���u�F�r�+û   u(�   �u�F���u�F�r�V��+��^�O���H���F��   �u�F���u�F�r�= }  s=   rAV��+��^������w��V��+��^������F3���t����V��+��^�   �����+|$(�|$a� �[ �8�2S��.�����"6����C��3��F��"q�*> ���#U�G"p�u��w&�]�n$��Restar�Ap/.Ox�!�`Themida!�TE!v���z�04-p1���5p�U��!�W�|���ń�`� ]���2
���	?�"0�y���A�tԋ���R��=��pD$�>�#�jE0�)h�t=�(�
%K�
HՅ�+��U����`�Z�� �3���E؍�@��~}c�t? ��3E��C��67�a&A��@F��|h�I�4 �E��
]ǅ"PP�
�ÈA�E��]u�'���Gd`u��$��[���7Tx�~�aKu�د�)GFJ#F�B�a���:����E�M��FF�>@)����40}��>�fmB�e�@J�e������°(3ۊ0��fr

9w��y3"a�?
f����
VAr
Fwo$Q]���9�}�r���v��� &���� �;U��Tx����8(�pp�Tp�� X5 �GIu��"�j�q��㰎�v7Qe6�܊&��AYk�Q��!���E%��	!AQĈ�� ߟLV=�ف�;a�yj{� ��$Z�n��: <U��z���b,���񚨀7�q� !eA�:^R\��4 g�9N[0v�Q=|�v;@Fu:	.�H��e�������T��S�
�)��q��v�D��0w"4���3u �A?�
����q�3����@E��J` b�R�M%�����Z��V0^��U��B2R'�չ#)�CA���K�֜��'�g���!@���"$0�Sqr ^.�W�o�T���U)؇��*Ԙ�� �����.�� ��*,nȆfh(�W���.S��0'��)2ϊ�[#fRZ�D�Md xBR��4np�w�qM� ��4���nB���O���?��v_\�
鐢�� ei�1�x7 ˋ��4�L�9��9�ސ���}���JO�T��	 g/R@&6:9`_��HsH��3��g�4܂�X�#�`��f��%[� ��* .�P�t>������p�r�v��Kg�������:�@C/����`�7�A&mXT) ��-E_����V�����0��8��p�vB���- �Ԡ�,4��"���>��̅�s��v�x�� t���dxb ���K%�=�>�NvE!6��������S ��=��q ���Tb��D)S�t��@��7� �y�<u��9/Hb =&-7@D����Ȏ�� R��7]�g�(q�3 �_�tӱF ȡ�!�uaQ1#�+�i�t�M)� �I۝��Š����r�:I�>�#R�d�U ��$*����]�c\� ��F��Q��0��� �
��Ro�K�����&�
�Ԁ��`��i���@h��`)�!pu� ����v�xW �[�� �$�(��{\`����0L�H�t��J� 8���h5���X�Mƕ[��-8Y� ��1����� +�%�J��� �=�U��0��]m���Oiw ��Z�j#]D���g�DKvS� k#�؃�����Cĺmϙ�D�h�
B@�yS�ա�Ɣ\Bx9 ���v �����c�� C�����:G��8-,9$�m�#�FX8LN��C�20,;�$5
��*����Xu���胐�fv���J��=���?��m�X1�� �I��Q%�� G bu� ��{���g��tVd�T�\< ~q-�F�1 =�]ӫ��P��t0�� �C3������@T�&�0���ƟJPԤجye:��u	4�n��W1�Y h7 �(p ����Q�C�0#o9d��$u��9Ô�G4�f�Z*m�@��ѽ9�L�TK��{�>.7�Ф�B�*-1�� ��Ͷc�� Ԭ��4n�Ͳ\$xs<%D�|`���$,�6j�0�����R@���� 4N�#�<0:cP��}�tK lv�e�A� ��!�ݍ� �HY��v�A�����-�/���.J�u��7o8���H��d�� ��;�B���z� P��r�������& ���Y��+�dt�X�r2�p<E��#�T&�!&Ɩ AS�ɊI�"����r`� ��F��a$)�+��ւ�)���CJ�q�M?`���&AO= 	<�c�X��P��_� �=乘��iR�4EI��@I-����oX���?�8�` A��y�Ұ �ʂ�G��!�,��Cq�,TL��m)�xYF	�q����@��.բ܀��(�8h�D�Z&X�<�/����j� u�VT`_���@�p
�ݤ�@6�� �l]M���a��F28da����U��\$Я���2#x2 �8�Z�I���Ά#��S�>R�! [z��G���J>`�5:�)=�(F���$ƅy���R���R�!qt�h 5@�C%��s�8?�{9�L"S(0��`�����:b�0ݸ�����% l�A0?T�G���&=�Pe��t&�Ы�v�3cC6ȳ�L�� ���1ߧ@ ���9e��$�B� Ih.T�V���A� ���d��#�6�p��<vY�W�ڐ�� -WѪ쒟�Dr�~ C��s@�Ƙ��m�d#PB�=e��8;��R�-6��F�� 1�5�VgrZ�Pw�\&!B�0�̄��5�.����pj��Q��I��`8���<��#�1�49Y����	*$,�| /�L!I�p��z#� l~$�G�ƛ&�� 87v@MU� �*12��
����<�v��$0�2������fX��8�$ʔ��<�J I�-��u�����=0�$�ö�8� ]\_( qZ֒v�94=R��>�ː �k�W�@y_VFn�����!��S���M:�5=�$(	E� ɒV�X�� 6N�E`�T@���ݦD 	ɫN�4p(���`��$Q?�BmM���:�� �����$�U��� 9��҅�H��j͟��\K] �H;�����;�)��u��@v��o�t�8��
�8���i��� 8����Xn(;�xu��Ѭ�I ��z2ٹ�����hx��ꩱ���<�[ �.�(�� �쾸|*	�TI������Y�~L ��PX/ rs:8����.�"�| ��� =������^ {���H(B�ϲ��8����Y`��:z w{�n�#�8A���T�<Ϲ��nȇ����&�N�i'v����0 �/�=]�l�0��Y�m0SZ@���+c Qo$ک� ��Z͉��� ޽H�f7_X��h ;h��~�;��;� G:�����3H.a�0�? S+��[{��J_H���/oK)���99�>��S'X@�(r��P�䂢 &X��ps
*c5�B�w���Pn(��5�������/C�y�.���!&�/�A����WP��P+�-e#X�nD q�b��:�� 0�y��Y�c��*@��$A�$��tk}���� �+��%��x�����ϠoB~�Y a�'͗���~� ����;{� Ys=ѩ��� ���(Ґ� ���7�� ��IA]l�wm �%"�=��0�@�Ϋ ��:�{��� �5C�ɕQx M�������(@�����$:��H�~��֑	����ؘ����=�B�B*L���"� >���Mz���@���� ��*Cv�� mU��H�֌Y(���� ��� ��ICxԌ�A ����1�� �z�R�������ބ8'����̤��� �7������ HC{ئQhM���8���{�>����?��x� |�kƥu 풩޻D��3UM@���� �� ���|�̊ �
Գ�"���Ӑ|����� 6y�����f����n� �Ψ��7� ����C��@�:����@d��(� ���*�F���0��n
�� ��7��N y������1 "����>C �Чw
ҿ �D���6������| ���FHo�X��"S��>�ę�7�@6u� .s�:���V4� k�^G� K��
dy�!M'AB��5�r��"ê<\ )y���-+چv!����1��' ��,�Ao�y_6��}h8� �*c�^0�gJ]���l�<�8ch�v� [��0X~E�@j�`Z��G�_�蹀:�<Ԋ��T'���i	��s�j��8`!*x�l\5/����� �F�mD������>�!h�mv'���֡ a=7^��p 5$մ�nz���g<�
C6�����������?�J�u�_7,@D�
(+��[�P�?�G�,6���K��@π�Cx����r���lCA���_�@������!j 1���3� ц� n��W�u�h|#: �����Dm�����G�9C���_@!�k@S�`Y�`7v�e��5�9�2�L|��q-�'���7o�� ��*�k�:�51"� �&�m��t�<� �PXN��=���[X�w����:#p afS�6}:�Xs+�	�wA�#T�BȲ36K]+���!�:��,�5B�r)�ػ��b@����@-�3
�7�L�vlH|`a�S�"�Ԉ�P�0_9Z������� �Uj����D�8}�T���>S'�,��
s�� '0~���G��˿��/R��;�����C"s ���>?�z���^!��x�3wD|@���?(C:����H���@	������� ߒ�z��`�X�4������ T@s�L4�ON�5��A����0L*� |R�|^0n9��_���ub�XO�,	.�(ZR����t�1͠�����0+�7;��	��w�
��v����3.��_�9�j7����^t�s!���9 l�[�>�/�O���Y�`t���s�8.=| �,�poLx��y  >����bu ��� ����^9O�d CS*�+���[�b Az�H��k� �*J��K$�� �-6\�;�0Q�����* +�D����XK� T�$q ٕ���C�
��0l� �i��I�	/��`L��XHT {P�74o�is8��� -��t�h/�iSrL�'C_Κ�t������@F|<G��$^@ľF�?28�vxҠ� ���� `�U�3,�JpH=F�HoB ��b������0�s���,ze�����r��@�����W.�P8F�mH��1:l�mrP�	B��dDH ��X����.������L�1�l�;��t�徤��tFu L��`Y�
J~B�܅��䐌�$@:t�5ȷ��ɑme�����4�Ĺ��p:i�/0�W�x������@bX6��L(���2T��sXk��)w �OT���U�b�l!�*�W'S;h#t0��r���d0߸�ؠ=��e$K P�,d>�&<��tF� �z��UbH��IҲ^��n�,��ro�j	h(5�`��]Jޞ3oW�T�8��������v?�
u���kP�JxAD��~r�������$� ���ltsLp$�����mC���DBg�m���G�tb@J"�H�3g7o;�#p��mB��C�f� m�W(��P�>/�z���C� e, :���:����X�m��3�,�c`�N�Fb���_I�W������v� r+}d�!ǘ!��?�����Y�������I�"< ���0�k8�=��r�=�is�ɚ�7wF���h-ITD,V �*1�e­x��j�2��:�D�����5�����hPs�1 0B�|( ��8�f�T/p# 4RNV��Se@X�|�D����`���RHKl@��76	�Eu���Q)����@�p��3��	B�v�@���Ow����%,�t{�yF�3V�ā�>�G��Hg0�PP`�"��h�4�(�@����>n?1�����$��dtFu} x���Qh����������Î�8���kRB� ƺv�\���S��
<i��}�)��: B�@R�3� D�Ϧ�?��}����)�Ze?N�ܫ5 H�
K�� �j�'��v]��ˈ�? �;#���a)�?,�XX�kP�l�.�Fy<D��3F��A�<�pը�7yZ�
P� J&)���� T�+�8�`G����pQ����r f� �Z�O�j���� /t5��;P�24�����p\E@�bg�,��LD�;�84�_��I=�-���H��p j8���g?}0d軃́,�a݁�ڄx��0He��\�ϸ�I��1<＂���z� {�ge@�v〸�M��:�0���7�Z��H�$��t0 �B�*�^�r�uĚ�� �=0'S�����hiz�,�L�v��D.�^FoH9
�7���|?�2� ���r4V߲Д���l`Խ���@H|.����6ݵ$4&�h@�5���(��h.LP�s%����������*�Ĺ26�](X`��œ ��(D�� �f~o�06�s����h�@;䪜�(�z�Za!8( ��+��1�m ��A�(p �02FX=�( q���� �; zȁ�#[0��ڌ��D� 4�Q�N�i~�t-�@r>�)�.��l�{?�y�����-H��t�7s�����Q@Xr�%�(,����s{�X+y �G�]�_Ke  ��F�X�����X�=���沀�G5�O���n��#������T���E �OS8s�`���G(�xJ����mG�Cœm�� �{`;� ��8���ζ��9`����q����[9�(�3� �AOI ��՜ �_�6���4�])��	���Ir8 �5"��bW {
�Ip�0k)���ꡆ�=��X7~��@H�h/��I�&�5���D ُ�k_�t'5dr��p�"	�e�AŰ�;a� @{O,PH�w'�r+$E��s`���|1��B2�T��d6q,�w��8W �`��\}m:�5tx<��|��ƌ9_P���ׯ��5,o0,��������~�| ���dj������VFn���~|����@�mf�K��>�w��z�W��@qo$gy����<p��BA�� �Fx>C��3>Ŀ@�;�䜜@��G ���D����>i���n^�|@�X/�Ѡ���, ����_�� tO$Q4m5�g���hjXAu��`�<�[0�3����b �,�����y���A����^�X ]KVL�A��OjI|^ 5�m�f��:�BOjh�@/8W��Q�ڜ���ju*|�{/�4%�fP�'`_6d�q�[��P�] �ޫ�*c�)'H�}�H��3f*,��@�h��s���Wu��%���h|�����7������`�@Er(�����l��+���3���?2�(QW`�G�v��0A��� ������f�<��O�N (gHDq`݅s��Ы9t�ρȌlu�+O��o�
�/�=�İE�*n o��.,"��SWB�� Q.�@J|�����[�&[G��%�iG��a���H���.U�/���]���;^g��SL�#=_�G=ݔI�rD6␴5���HL��|�+F��G�V��5��'�� �j"�e��,-�8%Hit�0��K/�������m �+6wK���H�p�&A� ٻz�lF��
�4��C6�>8�� ��d�����N�(�@�^%84�z:a/D u��婬��� ��.���Tu��`8�9���y%�?��{�sU�4��:c��Ls钡TéJ(��68[Tʤ�\�
@ ���@�/sD�� +4���"�ȿ�rܪ�&��>)��8��RM��}��I�7��`�2:���?��7�i�ru)���l�
���Z�nM�4�=��H�t�� l�5 ����0@N�<�|Y��1γ����w��@���~�3oP9��
�-����<\|��9z���r���$�G9��xT2���0�� �:6��@}�Ԙ��~��c xKS1H�l��6L��V��"n^	���z�&�\Xb'Ӹѽ��dG+�Dm�#0�?0���%j&d	�����1Qd��q���4C��8�����Ӊ�pd3PFxZC�%KL<��st+� ����� ��N��? si��R��$B2[Q��\㠜�;�D�3@f�G8"��5��E^tl�D��I�<��aR���!;/)�p'��R�%��A�8��������,��H���B(gq��4!Z�R�eP�����2�Bn`Ҳ%� @Ն(w�4 �������ɯ>�$�6T��!3�>�֖�O���_�D�����(�^��VP�H�J�`�ɳ��j�H�����q0�������!����D=`AKS�(B��$Ʈ���t�l �´�P�����8�|�4��B��8���(�O��H��-s�B�ݵ�rW�|�Ron��Xd��t�$OZ�����e��� ����06xJ�8h�
u�䤊h*d,� 86ꆩ�>��c9h� IB�l���I��!t(/�6��@L �=�@f��pf� ��@� ��A�7�hz��g�ǎD�K�4��ű_	<sܶ�&���K6�x{�H� 59CڄL=�ŖS(Ȕ�G"pWεb��:��Ӊ 8�J�G�_'D|�#�*s�@5lPߎ$K&)�U]�'�!E,3��ƃ����l�'7� e܎&��\�a�pr�	�uw! �eΑp���2s��/��X��3��oa�s�-�=��� �Abax�tp�u %)s�Q��#H lw��}g����+/�#>�h��z#0c�*�n:� �+[C���
�ٓ�����-;4 ��}y�Iuv�x����%V�`W	�[tp�B����e���r��Qڸ�7��<y�:$�x|�ha��$g���c�� 9�g��,%��M�����u�x�h�vyi�R����hט� ��P���T*����gD z6���@�wS�\;8���;��5���cұ#p�@0~�5���^�`|���tA9�� Z#�
��i��|�|��d�[E�Lr}�H i�%Z��� ��{ȸ��r�%�5�0�Z�$p�� ��|��,�p��XJ ��D\�<��R� )1+'`TMG �,���^���Uyc\��E�,�	�G4 ��;~���h��ԅ�B�W a���l��=MD�>�d��IC��D�q�x����\	9���� �g�K*#�+^���!d@7U(w婕`� '%S*aT-�(��.������:P#= �$�Js�1b��ëp:ֽ��|GC8\���@���AnNHSς	�h�&�pt0�A�2��8@|�/GcM0D��&�d�sV0���l����f\9O50��Z�FX�?|@jVIQ ����^R�9輮��B�:�&�/�r�.���}�8�N�PO�2�L�����bg~���J�>D�-�@�7�X;�5�(��F��mE��y<`i�m)���v@�	H�+�ܵ�D� �_�.�J�)T��n���~lo��ܢ@�ݭ@�3-�D p�Q��:�N���r�4o?�E��X�"���������0�[	Ub?�P(�Z��6��� �7I5|�� �N�>V,mZ�"
/����I� �:��{�\M���Z<� ���1S/���g�\@ �Mw�	�#E'	p��z( X��w3Jf�$H|*��Tv$� +���Ѳ�0[�7��_���UJ	�P����޴�>��; ��ҭJt<ր:�#r,�����q)��v˥ �m�*^�C%x��!� �N���f� �=jM��ز�p�?�P�Il�v��gu 	��Pwm�Q���z<���l�,H�kp�\74	�FP �l[��Z��B`�F�g�f��7� ��4HG���B�@ݡk-�1�m��;�#= L���O�1.�T�P��)*�s%��ٕDh������V�Ɂ��-"��ha�&@,ŀ-���x =d��� I`R����� ��$�8'��(� ��Y� ͦkQ�IO  �K�`ކ-��/;����ܠ{�{gMm@	�B����W9D��h@Լ95vӶX����U� I�h�ݔ���D�Q��<�\hi��+@�k. I�ښ��;�|J H�v��H�t�<�% <��e��H1�rį�0�?>L#sL��������n�����`�Ph�L�}��BKP�� 1E0JA��q���S�͆�y`}Ndq�K���f%�Bʄ@��sK�8�-)@�.:����iX�Pt�h�4�] 8{���S�����<*tu��3��<���s@ HPX��3�O/] �8w�x�� �ם�* 
�-��Z��4h����O���D�X`���/5_�9�4G= 7w4`ɀ��l {�y.)s1p΢w�
��v � �LO𙘀����-�/�^�����_sh����h{w�4����"�j0��O�$8�1ڰYWc����*�|�B��4�������6�� K<wl%:ڑls=����f�\�' 0�"姂y�	;�*��tFn�3�9�܀Ʋs�S�����t���@���5��_���rA�/�#����<V����~w����(LE�  8_(�hx
���������� ��crjsm�)��ԈPZ���_#0rE�Є���lf��x�� �*�%),��d!�!��* Mi8�� �A�
�2�ɫ�tw��.����r���/*���@d=��t'������z(��z��C�$&G��qt��5ȯ`"��P@?6�;����P��\�������~/m!8�j-��g`��^F<O���w+�����>�e�}��Ԃ���< O��HB�~��,�o1� V�R�)p+���&�1�?�*<��-E���g0ڪ�f<5�i�Ȁt� �	d���i\a��14��d�$^F@ ��j���,.���)Ҵ�� Ckp�?GP�+In�]�8��i��-C(�����A�� g�w�*K����%ҵ��1X(8�z��%~���)��Bn�^��i� ��jn 3�������8������K���!o�$/)��mw�_�. yݔ�џ�0��I �P��L��E����x�������i�-���yTy=H��ks�޶� �u� ��"M���(� ����/m�P�(!�J8<H���}���!�Q����,��S.�(�\ �ZV���R����]�Ѝ�,.�!O,` �Sy��E�,��2��J��$*�P�� ܢ�E��Jkh�S�p#*�db��1@�E�C`t�(v5p�L���2b%��Q�A�=� �_f��g��~7`�^������ Y���r�v ���NU�s���J��`����я�@���zӽX��.7!��,08@��F��6�@�^�,n<L�	&	|?kA�LXV tu$o�/���S�̬t�BX�u�����!@�"�z���������@��@�(�%D���p	�\'�*q�<�n��ܞDo{D���R��8u	��4�^,���X�� ��.��7�� ���n(�}8H,|?��5��PT���>�'B��^F@ =�����M��J��T=��- \2<��8��7o�^<��	
s��R����X{�Y�B��HLr��d�� ^ă�N+aedA���7?��R �o_
w�E�*6+~��t[(R�'V�Ө�"X9@@����A�-�h7��sZ���'ꀩ�����%���L �]�Z�缠~X|	һh*y��v B�ؘn �_F��l �Q"��>馨�pfĄ��0��I� � �20nC8�a���ٶ����,	s�:؈��i���"�'
*�帘� ���Ӓ�A)E$�mbvW`6�'�#��ۆ%�m��!� �l���[I��t�"v �qdx��&KDG�s���0��&�r��)T���'�[5DD�c/���s��3p勢�%)��� >�LB=�^.ػ(����s�Z�	AR��5X����/ �k��En�.�è��p*s�s��(ڜ�����	{��X@DrĮ�W,��(p|��繴&�tJ�7��P08�@�'�X0N����I[Т}���Y?��P��lC��H�H�_5whd@Y"c��"��)s�%���\b��%�D�Z�кG�^[g<`m�
ƀ[��?@5o���]ΰ�T�_s!�ҳz�:l�D��ot���@��6��BK�� �sZ� hmP� ��;�CUʱ�����@�{�5�x��?�nX�D�)n��#�R��! �J�|t>ٔ}I�9���1 i\��uܨ �Q��� 12 ò	:D���+Y�ڌ q�ҔA�ۅ��\�t-�����ODU�QGp�ɤ�|�m��k���<�K� JOU]j�_�q.�e��	��h/� s=���Ԍ�Xc�ޯ8�4lk|��Å��j�h(Ԓ�S�(���[X�^ ��/9+��t)-�n�@�o��+�l@D:��"- }��t.�2��c���Z�����J<�6ۈ�	֬��0'B4�s�u���˷%���$2�,9�l?�5��H#�Ĳlh�ȩ�'�� 5�̩���؈%��I,��t���"�m�D*�����P������W*Tp���5�.@�-�)�S@ )��Ϩ0I��\,	C�l��H䓜-�[�h]		ҁ�p=^�\��U�R7� ��1:�oq�z��b���5 ��(8�f�Y�]�9�> y1��9<�#�����	�w� 1�CJ���lB	@�7c��|���#/󀵙�(���[���!�(��1�M��_�P�E�9ɜ�h�1��F�d۶E�@t%ĩ�C
Č]��G�\ƀR��P�1 e1�~�Ӎ5
ٍRģaA�!"rW@u�b��Il�6�@O�@K�b�(�,!�Τ�)�&\�sx -p1d% ���FD�ˉb�H�$W�I~Dė�(��X bWQ��23�Q�����0�mY �0��F	[&��9T%�?bs)�����$\L�%;�@��@P����$�Ib�V�F
� 	�3�` �&9:0�X�P���S�` x�Tj�=@�d�� G���A�!�1�&
��aHDj�D\C�w�i@kb1d"r I�U��܎H�E�i�p<� g� 0Sά�:��8�M�D��j�2�" �����7��Ƹ�� �6
��PWQ�砇Y�'k ����`��ڡ����5?�(���[}�KS�t� j��&5ژČ(�ҙ��@~Bl�LP{� _�GC6�JB0�� ������C�栞p>{�+�+C����
Ѿ�p �D|X+B�.h�U��Z�R@�� e΢1��m�(�R���,�0�JE<+� L�m��U<�/'� #��1xj!k�Й�8Qfˉ ��?y8 �+��E6�K��!�������L	�ķ��RPړ0��p;�:$�+�@����ؼ�r\��h�/����@ x+}-�J]5=K��pW A x�d��V�r
�Bб�@vǼ w�8R��} T5]����[r���#�
�k��B�lZH p;}�h`�>�ƨ1o�S}���L��uGB@����(9�
�0k�� ]_�<-� �ٝ��D�i ժB�Q�� ���-�#�G8������Y����>���f�:'`���u+�t?\� ���EHAH��X� ��Q�Ӏ�T>����@C�k�xYB���s�I���|H��jV xw��q��(� �e�,�X �|����(C���@�cmsA+�] 3,�y��L"x7�±Sv4�0��@��q�-����Q/Tn��@Y�:�k�,�m�"C@0�iL���1A4p�3�|�c�n���`%�K��<� o�BP~�c{H�H�i�mҰE��ԓ2�Hl�T������� �IٔxBT�@�+מh�(.��4DG}Bog(������#,�	[� �q!B��03��S�� ���$"0W��G 3�+������2��x��y�Ň3 �P�%_ �W,h�^[�\FD]�xǀ����1�p�w �`+߸��$�F`���Q83��� �x�X(A|�FOG,��L���p$��H��(�d����8��&�1���0�@�b?!��0f�`+��@�^���ë�T������~Γ\TE[��Dhh��#o��1+؀[��'�[3��r@�d	L�E4/�9IdW��R���[ ��� ���#�_j�*Bs	Puc<r	a��[1��8���$�Q�ʥ�����Q���*`�X�M�� j�y�0c�i ��~E� Bv����J�Y��h�m���!fK�Tc��鬲0��@l� F�j���B�:�r
�K���0`�p�e��P�|�O*������u����1`ا ��.-٘H*��$��}Pϩ�3������H�H��K��#��I�X��&' ��h�tK}3B�t�;����٘���D��k���BL��� c�|�(�#Y=��P���| A!��BT2��x-*}S��qh �D��x\Z� �x< `�ì3��<�q�����J� }�?�j��Tz �vC|� ۯ���5P���n�|B~D�-�+��}�r0t�v�U��$,�@�%�����X'*6��n �;�}�������&�l��D�Z�gk	�.Bz(���R����؁0�/��L	�p/�Ji��\~:c�)��@�3x��4hz0�H�KLT�+�B���W~_����R���@Zl=��+��	E�H�"4�Qb�`���D� �r�gB(I	k��܈��> Hdc�������J�@ PЊh[��,�1$d�%���C��C���zB`FXW�� �Q(�{<�\ 1��h^�V���хu���� �3K�eCh�<X� �, �_.d/4�;+�Wr j��*�RBg`0��K�H�d�:y��F�D$�>�Ѭ�3`D������*�P�lr����A�F�0@EXAܮ[RD����d��&���	R`a�(m��ڙX]{3NKKT�&��&�i$d@�q�,��l����|{��Db��X.C��V-5T�d�W:�>�d�������pЈA�15=�3���	�X� �:�2�$� x��7 ��^���,�5�Bfo���J��Z�.EHBB�	4���"�d�;:�j��÷ �zD�Q6�%� �٢i�}DlNؿg5(B������ j�+\������E����5�P��,0�˼6� �|�Ӄ�I,]�'��h�M$aH@���]�hz�h�V��p�rs�0�� �+�)e�z�dwPU�H%� ���V�?��%�����j���z�t��Ɨ�̉>�L�ki�$H�����`<b�+iP�8��:X��1����ดh�k۱o.�p���B(�t�	��5$�ց�D� k��tZ��������pA(6?�t�B5�PH��Ia�:}�;kE��r� �tC}|�]h�l1�B��	h�� P��zL�@&5l	��� (��ք�P�;(�ԨD6|�yB��: Q&�����[��@� ��/B�?��\� �����?����A�`)�m��s�r���?I��^
:����+/���
 �j��*�ܫ�,�(
)��|I�$(�Dv�\P���� a����\72 ]ǂlBF"����&p@P>��x�`��aw���Oy�D0��n�s�c�<����ړ��{�j���">� �}��F(BP6��3̨�`E7J��;�i�j���*�t�ڑ�-��l�@��/��Q�ǤH�����5�j��(�9B��dT�	"�=Z�H_� ���AJPT
��w:��\*��B\x�S�F�1�M@�EH���,�L� P�k�6�Aq%�i\\�<��ÜV �+�P�O7���(t�xȼL�y'B��0�k>�*�x=�4����w\�x:H ����]�:����'Wk<q�`*{٠5��}!Pl����㒳b,�x6���	�BZ���iTw���]�= 9��6z�� �C���'�����%K��`Z���u+B$��
�~��V.�h����ov'A�(1 j	m�b�Lu�c1P~��<����{ՅD ��k�ǲ#u��p��(a "�[�5�ɴ0�?r��Ă����p�;,���(NdB��ؼ�l��,���b`��v �Z�%T��AH� '�����Y&)��q+���b�.������ķXV
s�۴���X�{�r!xyLM8����uC��yi�$a+_ Ŧ�rt�\&P�� 0��R���' �MT4�%�����p���XH1���� ig���B�	�`<�e�E5�ԁ� ��� �CW2jo��%"�V�$ ;(���|���� <�I(�,���:�A���u;�p��n�جe���"�`L�D�O!TQU�xԌ=�S@��(tc� Pr�� ���� xO�9=��X]�@ АdrB�6 ��0�,8g�w�!&/�٢* `6D`Ƅ���� ��BV|�`,3�.��qF �ګԄZu-Ӓ �W3�H`�8��+��X�<"P\	h�+�ͭV�BF� �qGUh*3�Zn<�����(��這F;n� k��YQ��I(,�r���� �59TlܑaZ��G�R$��tv�h�k�8�n�`I�:�>�2�Bg
�.� m�Lڔ�d���ARvW�zD,mn���8� ��/{ *E,�ԓ�!y3����0�d�G�P��R;J�ȜQ0�ˑ�|}� ��Â�p�iC�j��u.t�����@L��`�D@\{���axc0;���� ̦����$�׸�<�D,��x���ȳ{���ޘ��`d0G(*,��b�h��]/������K 늸�J�ۑl@��,���B�l�����*�=�X &�	K�tC�D�0���!���܁ctH�y���KƤ�0�_kv���ԋX��\əH$:�R, ݺ_� �D�j��JZ���P�����ti���k} ���k� �{��nC����G�H��kRȄg`��,�_b}�PI	t�0:( 1�VWn�QT�"c���k�2��ҷ� 0/��)��Z�G�J�	8�.\���AN [��X���kGh/����	��4(x!�� '$:xB0���`�6�i��k`��5'����ÅyH؈K0&���l����3�x����9ڈ4di� 0N�4WBrD���J 2��Ӵ� ڕ݅�%A�(���P:�@�W�'�p�ק���L� }PT,P�Z,���,
Ҷ8� ~��4�#���8a��B0��Ѱx�P�Ny��7�@�=�+j�1o�$R�d�����8 ^�1,*������uE�B0��Z��K��r� ��Jcӳ ��g�6��\Q;�j
����H��l�B>@\�_5q�ၔ�j/�8����4� DP��!�Wc��L���@{O�a<ˋ���L�v��h Pz^$� j�*�,y�C�<���ٝt*��+�mo@kc�O�Pu����]8a�ň�+�8�PDP�^��p��x҄�\ �ܗ��`\��q:0��+���PC�SU����B|�\�)D|�^�k���yp-� ��<�V����u��͐62�p'.�3�XC0@���;�4����9��-�pV�C�z�%�� `)f�6� d Bn���=���>�X�����9����� Khx��ZC_�]h�X�u ���ڟ6�`
�&ʬ�J�V�� �j��(#;y�$� 3K]0dj#<��̊%�K�P-;��� ����ޟ%BO��� [���\���X�����  �֍���z:���䔰��tc�<`t�1���du�3Ј\hi�x@���9x�n4gy$a�p�"0����\@��i��?B���\(���H9�8k�D�HjU +���~D�E��*@���7B�H�-�x+Kl�k�,� �4`��~��
s�O�8�΃���A�+ ߜY���N~)�blo ��KB�j���X�4�􃓭�@���v�X;�B��X	kL�^����O�8?�#�VC�:��>�
[s�-�+P$�F�PB�cxe���"k�9U�z1�u���e0 �^UK$t�3�"� ��Aʧ����ip�B� ��0�X��|���Ņ��`�K'��k��*�<0pal�;(|�J�*z�0�xٜ� ��:�+��B{q����!�G�܀ڜO�)�s�zp���3���$4$� 9Q�(N	=?��4Bs{(���w�� t�g�%x�������� ��9�{�6��l��7�TN`^�Ą�<�p;�T�<p���1��K��:D��ZqXB�0��5���y �7�P��pϡ:XDlZ1�րY^|��|�Q�}��r,�o�d�"�r�F8z���� �"���>}k .ړ�ث}rt��x�����B-!��0e���h� �>��ɨH�R�� �|���LZX Ȼd
�>�.�F� �-�؄^� Cwr��T�:@��0�Y��ҁA�}�	+!��4�S���n1��ek5ȘLA8��^  |�� �L(�K��rp��e�<�2`�TP(�0���F,�8Q����r^��ze�9p4���_w���:�_� ژ`�,���N��Գ�6�g�����O$,���TWːK�`��G�T�� �r���M�*I���p	�B'�v</�t�����h	�uE �B R�Д%�� ��jޑ��^X� �ܥә�K�!\y��:`���w���XTVğA��&�8	���ͪ���2~�8lA�1`�B&����`�>��L"����펀��~Q�Ȋ$�	'禷,͘B�`���5�H� ���Zs�	B�?'H<��%�1�H��]I�Q�*0|�?��B7PД� �ڑa���,i�ւ�T i����?2�q��$�;g `�
(C_6$X������d'��<D�>5������:T(�}�������yB?��Z�������$t��xB���Ę���w1 k���E*�����/BL>ipxJ��s"�xన�-��b�Z��� �pc���'1U�@�"d?z��Q�as9"��pdA@���8O����@�fZ[�w�X
��`T@@,G8��PJ 9�'�<�:a�W�j����G�i��3߁YoBW���|��w��@�=3�ߨ��ܨ ��t����0xBp����˱d�0D���x�1R�����������l�#�Ҹ��V��7����[@�D��B�$�ј�:��'aB�8*�kg :�# 7��k�����O��Jq��{1�ichZ6h/��B�\`����D+>d0W�\�އ�e�Z?��������.J���PA��`��~��@2j����?���C� &HVX�{D�:����xP� ���Q0�>�	��
��D(�H��ɂ����0]��z�$NP|o q�X�A�8@Ŷk�/�c8'���HM�u@���X���;�1`�]z}���B6� P��(@��3ˏN�l�ޘ�^�(JBZ<?tt�	�#��\g�`��|���H3T[�tb��/��o���n̩b�8�mlQ�ft�m�p�<�#���h�֊��X��? ���ꉷ+� a��Z�K	�%�� �34�ok�)�Z�.9���O���B"ު��/������J4��h~ �Q���-H���+���{��$d䠨G^�ȁӸ-�p��,�+B{�N��d�; ���(?�=�4Z;�E$F ��}�:���L��/�`(.��-�T�+�T͢ȏ�l�� �����%4��GP0%qc)�#�VL����~��;,���%jH����<L3��q:j0�3ۅZyC\젳r�*[	�mӨ��=���cQ���P<w'�܁p�B��=�G��F�wi���D�|�l�@ޭa���d�G('��� r��0h�@����s,�$�G"[�_&z�O���Ѱ ��{}����q#��<z�r�2���� �WPX1������0P�p �/B����Q�cT��h� <��B��@<��HX� �����#U���D�Ґ�	XS�v� ��(�Q�0i��K���f�-�>�(F�N˩�M4�<�N��j.(B��P �g�Lʌ���k5���[D � ٠�\i�d�L3�_�p��0 �?y��@~8	��tU� i��bkB`2�ĉ(!uh�d�p)�C ڟ��o��_��,6s;Å�ɖ �LL��X�ژ� ;-�jX�,|	��(�L��zcUO��@Z�!���%<@�#"<{A|B��X�%��K�@���ڔ�|�kgi��DB#DlN�z����Ze�x%ځ��+���2y��nC��!(`��/N����rP�]Q<�ȓxR�� ��^��G���E�4,K�(0�Z�I1���\�`�B�t��D�J�{d�ڌIL�HlL����O}��Bf8n��/�@�w�/[��B4ھ	������	�ҭ�Ĉ8Qo�i��+�t��)�,S�x9BXT��L�%�E pGbq�~�(��42�x0B�Xj�*��Ym����J� �^�� E�i���x � �L��*��iS9�-'z0D5k	;{�+�Ly�h/�d�)��'D��(���x.�٨��DֱI<p�\jX�Bw�TR���@��q ��J`^P.u+�̎���� |A�niU~�}��+�vʆ�
'V,����X@pS�0���.�.T���	t+I����;�q�xC��$��0���
 8P��/�5OB�r�r D��B ��� @�b�$IT�uBT�~Ă
6�@4� Brڝ�YC�����u�[�ӣ4�� ���XT�;����؄P�A��S0�Y�u1ܥI�d��:�'��H�
��a,D��4l����h�p�P~_�2���ҍ�0|� [u�'|)��`B��@��� q?8y��e��9�ʤ	���$ [�HvP���Z5�x� �K�FP,,��IoB�'p�yb�x:Iw�x���|�>L�d�x���9�F�5����lx�:w��+��-��@T8�l$�-Y kq���w��@e"P������Q�l��W$ @?��/5ZP�Bx���p���H�F�G<BdI���W2۴�:�%56��N�+��)�4��K�8慝8$�b�=~���\H���X�V���[�*��H'u�hř�����V (������DA�˰���LwX�PX�,����&��(�2�I �`��Rl|\�J �Z��A���ye�;��%X*�.��D��0]r�� ��ٛ�E�!}j�1��9�����H��\@%A'q��T�*��1
�%��4�0�pb혩�C� H�>�i<�� ��Gy���E�0C�Q���0>�`*�y���0�p��}�j� \����� �����*��|�:���G0�¤�=�!����d�Pr�`j�h��( !X�Dw��P`��iq� .�ٜ�;����Af�%W���z>�j -�n�K�� i�sU�Y� tR|,�*�a����}��c�oj�����������l�3��iꨀ٘��jr$��"FYpD�A:�@ګW0/@�~qp|Q�����L4A5��@�� lF(�+�H� b�d����يz�X�i[�>�)l�H����z#p.��Q�����(i�$  A�t��1�Z��O���[���|gNI��i� 0�l��|�B�\D���q� W!þ�)|E�01�H��сJ�wAe����(/ I2|;�􇋵��������� ��'��d+���2Ѻy������\����*��x<Β (�f,�C�H%~ )�*��MY���4J`��I�6P��� ӧ.H�]�DㄎT��4�8����*J��q���>�D@`y��`��Ҵ���8�0�@��਑\NR	p@|rtB:����+W�;�6�lAO��İ	�k ����Wz�,J|��	)� ����Y�Dxq9V�j�)�b���AWT���m ��)�������׉ N���=z��qA��P �"]U(:EL=� ْ�?d�G�>�$ � �:�o�zҁ���Y���L���&p {�9�<��Y�tBȐ�o�{A�-���@�v�	�ڽ�����l��PN\FcH���a����B×
3�$>a �Oz��� r�����a](��F�Aߨ�o��Y��hH��O�Ւzɀ�A'5�I��S��` 4<H~;��ժ�{SHT(���0�A(���� v� ]sR����ay0�� �P�������` �[տNvA��#��YazP�8�� L�0��(b�H+>�������� ��e~�١�p�������-���R�P@�c��� W`���k !����d��a��P"��s0��H&�{#w�գ�@ �.׭�M˅�)ƀ�fr��~����i�f�p+����qý �r��_1�0~0A�U� 9�ʘka䲯��.p�

f�X1�
j�A�m�����&�2����������>2im����~�I`�� ���*�Ð=���$`�.��x-�~y1F����%\��A]}�X��&ƠTsy?���beB ���g+��>� �9*`�A�� a�~�����C	�D��:P��m���~��̏$wHT�����P����@�i*_ܰ��Y�Z�����c� ��`H�{�� �'��Z�7��0�)�a�*ei V_"ֻ�����p���+�� ��.�h�G@�v����1�����%��N|������Z�b'���aR(�����A #[8��&� v�\��}��[q�V@�o!8�%�Z���0��e���P��i���lz���0@��.�#\`
���� ��Ǟy�x_
6��(�p���l��{��&Ę����.p�z�X)��A�i��#��y�s�*����.�x��Q��� ����`�� ���(�Ah��%Ѡgu0ĝ�Vy`�P�������,(�0A�ʡ������.{t(L>\�I �4)0,]#Y�Y�q��%ձɌ������U��b9	�����P[Y� m�%�*q���Zs}'t�G�$�f�� ��q)�HC���M!xP(i��ܣ��� ��8�&��������4�L�4�𘴋0�@S�i��y X%���J�p"������|W>�심T���_� ���[�i�8�&��P 苣�@��� �g���$��� `	���2��rό��@�\ �m���h^8�e SWM&�U�"�b os�����`�g
�L���_~=���
� �i�ͼ���t�X
R�����$��(!�
���B�႔h��_�^��~��X�NRӠ���!# �֖�]�~Y���љ*��!C��L8��!��2t&�&�p�)��>�V�4 ����H��I��iYa-�'
 <�~#% T:\�x���=0-G���A����D������(H������jp�`���Pı%���4���.��t���ٶ����`�a�G�D��%@W��u��#}[^��A�Zlв+�q�v�X�XW#X�$�. �R�����|\A�� ҂� �7)��r����� ��T�q��p*c!�"xV����&���{���P�����S�ɤ0DW �#�C]L�<��{�~J�����sc랎T��,A�� �E*do�H/|hP��ۋ4 @��2�5M�!e  
&*׀�<��S0$�h`��fB(a�� ��%,AP�� �=��J�p0���%%�  �n��o� >����rս�t���y��_˅nh�f���$|b~�hjSʎ[��

�����{��} w�)+��&� �Q�h'Ţ`��S8���R[��~36�x����=Y1`РV��3�i�ySX�K�����Vܣ�����Y�P.e�0H~0QĀ��� 6�m Ds�0`�oʒ�Y����\C�˧����h�˰@�S	(Ð��� ���׋� �c�l ����hQ�����ȸ)��dhX����Tj�*j��XD�pZ
 ���ctF�*�$w �X�V=�0uH"r���sx'�P �T�M �4n������ ZG��V�	���`Ǐ_+iu� PU�� m/
�~�p��cy��e������囀8���}�Ã��¢�K�	`��#8�s�gQؠ�~�SZ�T0�VP��'M������	+w�ХxS�؆� j��D^��� iȴ �0��0(�\L$�P��~� ^�ǂ��� ���f;�Q]�ty��&��H�\,��`.Y���m�R�D����ٹ����ꘓ�_�*�pІ ^Ղ�2V|���G)43�`��c�P�v��qItf��~e1�f9����������z��S[���d0� ����q[�� �\������TІ;�B#Zq���q�ತ��!���Ўs(X^�����	I��.���d�X��7� Z�]�a����Б�pdD=�Ob�kP�RZ���֎�-B�4�@��PĐR�(�!� �P�X�X�\��$��T����6�V�t ��<�s�C`�N���`H{���mp#]O�0⎍�����l�A�X�%��tZb|���ЎWت܀,�"�n[���U�}�c���f�B!E	&��p� ��d =��۾���7Ӓ�@�IN��@����ޥ�:'x �(£�q�����x� &Ř��ga	��Zt��{'�Q(�@����"����=S��@������~�J����2 x�Rh����~��_�����T#[�Rf� ��-n�8�av��B��(�ǀ�	Q�i	)��� � �+��KsEX���
�줵��� �&�(��5�O����!�~Y��P��Gİ�D�ڬ	�P�(�/��BQ�'L�',ꀦ<֛��vƙ��T��`�9h��������tr4 S��u���m�}\+�1.�,��^�'�2<X�x�� d�O=I4��
:O�$d�����`WP�~��hc�X��*�@����}!#�3SZ�@�W��C��'��<U5씈�ԃ~}h-�,`� �fH냀p����@$WhN@_*��\��c)4$�����^wX1���W�E���Y��^ ��s��U<M����_:�������gO~�:� �8U��j�X�3Ib]�7����W�L�"���ψ -�:�@[1u����dr:<:�jb�8� Q�c�R�(�f(��3Rs��`�XV�	ķp�\��P��h*�0��D4,�T��)�X�vo�1SU#��[��^��:��@�B聀�	57N?)�Q�	�l@Ar)oL�DBYZA5���������Vh6����$��IAUh���d��_�Q��C

	�^��jI,4���wL�� WIƮ��(H[?����p�4]P���4��s#f(�H>�$��^V�3������怊��^Y��8֐P`��X@5}j�� �n9��.LM�>���U����2dU fY��h�T�*��u�I��9�:�0�h@W�5<$�@��P�t|X���"W��c׃4��-�|3Ax2�5����5�	�RI�Z��1��7�~'����\���M�  Sh��_���/
�^�0r~jG��xi>Ƌ���3��� o!%)�S�9�R�8���i���{�V�n����Ȏ�G���ZRTZxW �am�'!��&����NW<gގ^b�haM߁&�݀���ò?(��gs��D8�h j7��&Z-d$j6>���P�	Y�\��t���;=���׳ϝ��O��[Q����S��q۪X��GT�<�&Z�)4���Q$� �HSt�$�	[R�]�r��)�-	}�C:7�~	1�;ҭHٌ�R��o�r�:��,�L�����k�@6�Y���1�Yd���|��)�H��[��*|YF����.1΋E��1#mݚ��4k7��՘:f܎:(h��ĲW��'%3�1�\!�_�b���9㨿��Fɋ��_��$��\ܴ�R��#Ih����ꏚ���^"��5�&0�OS �=�$�
���Z�����C��3�ۋ[�E�`z
)�2"g<Oq�tc�U��8�@���k� )�Y���ݰ�h[7��DL��<TM�����D�OHF %��qe0dL�y��SLB���I���y>���1�r���!=�X,)�* zZ�n���(m�駓U
��h,�J?j==Yy�v&2�E^@d��ұ���!.��{�:BH�T��,�i��LW9�����#�$�\��hUK�c�*tgn��и���W	B��@S�G ��5	=d�YA���x�iR�!�
�s�G hEK`�.r)Y,��������0��YN{A&"r˷�����P�+ ]���p����O|��0,�����Q���l�Ϗw"`v棊�E��YV@��Z�f�g(M���-Ә"��z�%��  ��jBkh2`���]E�^�	)��&� U�j kQ�Ձů ƀ�]顙�Y��!u�)�D,t!�ba��� �E� �FH��6��%
\PTX�I����$$��d�E�<=PDZ1�ar	�h%�(�V��c�]��v�JL�rՕKLB1	�hc,���"��*�� ��eN3h�M��+�Y���� @���%��}� ^���T���}d`5��zX:�,O,љ�<2`���ӿ�V�{a���bs�W��cZ;��&�3q��B�U�]PLR�#�Z*)�
DXhX鱏A3�]&#)�h	 �t�1�ΰ�hNi����@Q9v�=U��"3�\_^���FI�L>�ߔs}H�� �*���V��k��.-lI�v�ʑ�M������@Q!H�LQ������U�7��_C��L`�M�0k�һ�y�H�@.)�X�YR�JR �����Z��3Lf��o�j!�@�Tg�}J��F4/:C��B�	N_1�F�)�X�	�JZ�^c1� q�~�-�&�=���%���^� ��%��� �1��4VMF�@ �".^X�371h5�5|vX�RT{'P��6t~Sh��B�hDB%E	�)0MY��HR��$�D�����vja)� ���ZDm��Z&�����̷��餿v@̀r�ʾ �p��>�O�!�Z�'#�f��]v��qh]/>ZX����~A���&�H�4p����?]o��]��h�YK0���8��N�@�ƥ-(()���Y77v)�r��{'
0��b���Vh�r�X ^Q��#~:1�Y��q?@��r�g��OE@&qW�i1$�Yh��doUy�S
*���=B89j�
h�T�d����,k�\	_#;��s���f�;i���H�>2)}�6wN8F�%�l�D��e�($�3F��`�E.��=z�[ f�e鬼(+=�7A90�%IX1���\Q�VQ�k#=T���c�L9X�H��_8�|ׁ��E"�4`>�d�����R�0�q^Y���2&A �^\F�)����c}WTJ �Y@�
!(�S$�]
��l_��,KWbh�,EK��cSh��d܋��Q^�{������W��g`�|L
N�=��&F0h{-~��{n+D@�����J�C\E���.ys�	�A��p�2�����"iWA���6R2�Vŉ�pD,�	�8� 3�oF	N����"v|Ӈ���v%O3�1�vΓ����.��F<�¥����E�c�6��i�T��B��T	[�,��==/&;'�&��U,}O3���A@t-Pb�ŝ��a2@Y%)�2w�g�dh�l����p��Ѭ$��
[�>�� ɀ�{]1��]#T��}��s�!cD���h0ޫ����� T�$�)�|-{j�v�{��3P0�qI������b��H\� �O,�9h�[2 �e3���P���-Nt<�
�>�XS�K,�g�E��q<�2��S	3���u
�hCV���-�״O� �#pu��
c��B�� 	�Y��B�Cd[��,V논@�؊\h� ���y���GK1������Z���μ��3�l1\f�!������0�HX�����1�･9��b8K��뒇��-�3 >[����X��@�(�/���Y.(��0��"�����D��[	 ��PQ9��-�i�l`�3������ ~8�v/��ARG҆� �� r��
~���GN�� �"ډ��Y,�j{��23,���6�y)�۟����^@�X�ׁ�6�Q*���L�*��4LI.N|iSU��Yl�W
�3K�(  ����[��I�Q[���=�&� ��w��&�yMaY��2�����q�	R��#�{A���:�q��&Q��W,5�D��5�b�PߵBU�o����3����g����f9�v�J/:��(<AC(���L�	����Z%tŬ,O��0� U��� ��K�$ʼ�`�MBS���N�`j6V���I�[2�fQPR��9ꏉ�n���������R��3X_���i���T���V�S^-�Wv5���j�BGOh��oUk_���� X;"�M��o�j�*�Ř�_Jh&�����2�L9Ls>Oq��������(��3Y"h@*0��b��f�	�Ҷ/p˷�V�.��Z�#� T�w�fY�ӵ^��ݏ�G�V�P�R\�E��߅1U��@�� �iT�X����V7�e��m�s.����I-SV~�� ���<�]��X��1����IJ���p�LP���;Ac��Ѹ	+a؃�B�iBW�Y��b��^��# 5=(v	Ø�'�Cc��?wN�INQ	t2gB�Fm |E�#�j�Պ�H<	�_����H��c�
� �4"��L)ss`��	2����$�C��$�
w�R���3�\$��	D�h�G<2��P����@�+I1X����x<��lB	O.��[U�1!(��,>�B!�m��v�3����h���Oz �U�A�SMQDɒ\P�؎��uʤ?�g>�Ғ����h.d"�`S���[� �*�ˀ��Q��,[
��hnKB1`��$�ƟC ����Q�.(k�&sq�J{�@'���� �h	{�� ��n��y��/=:�|>J�uO`6�B,�I)�7�mcP��ݕ�b�8�yc�bKHЦ�ԝ1�[W���`�r�q�)��ʠ�-�H�Lgd)���c����X���҅]KA-u��6�&(�&��|��`u�y.D)U����Ph�;��+U��.A��(��)�;�SEmT^��+a�i��K�Z�(4��վa�_���;+\%��0�=\	�:��H1�X��f��!�fY���n����X����� -�z;$ª�F� �ځ�,~�;�8�8�=�������P
hk����iY'8�J"AՄl]�;J\(�S�f����h3F���'���S_`cպ��HwF�I�<��/��@�}/�����`W�Q0�e0�tW\i��"J#}N� �($`�	�%�c�p��+-��{4)w�X���9.c�4�������[�����@i=qT���݃�Pj�s ��� �p1�])�Z�" ����X��/ fh'铅̸�y'�c,�(�YQ�a���S� ����j�9��	�]Xy��j!7�E˥�î�P��[9�h�՝��I�W*�����(Ն�A%�DX�vKP���;�Qb��,�T8��K���B4	�
;hk3`t���Qͨh6;V*������Q�̀PT�R��
<c�%���5'L��0�D0/]�����<��X鍆!����u��bh�h��ܶN ����J��cyل_P�A�{�X��3iB��n̖ Ƽ,����ʀ%-f����� ��t���[��H�Bn��.Zsi�G�i
�=w]�F<��2�yT����8h�t7�����p{�C*}9�Q��z�J��1����Z��X0J��wLP�Ǵ�)���,G�����bN�V)�R"�\�eo�ps-@�3���������ݷ4�	��R���b��C�4�$�H���f����WZ,�MAH��"�B�QV����K4c񌧳��q�K%�UĶv].:Eai=e�-v9��A���aE�C����+�.0�^�[�qu��ؠy2фF�0x'��z)����ZSܓ�_����P�ST[hHg��5
���h�B#/fXDF̚���rs-�kL|����&���HI9_Y�I�KWT@�&#�
2�`j�Ʈ�o	#���2w^���GHyN	Uj����Y&��L�K��Y���m�� ���T{����ۍ����]10K3���Z�"���]1� e<|����@�h,wVi �DB`��rZP�u}�F�ޓ�ܩ�-��b�S[t>��c�,��	���9�!�%���_;�(�:��b�@Y(0P`e�S��������<�O��'_��RO0^��IK;f>�u=�A����c <})���(�PAĭ�=�W�0!~ 3OS���u�)�[z�4r��s�P�ًb��`�rM4��} 7Lo�>)˽���i@޴9Q�Av���?&!iP.x��OW�v���z���#`������[S�,���t��@z����p{e�1��z@��� �R���ڢ­bB�������+\b� )QN#]'��@*�r	���U��.�Sǽz �e����\�0��h$�E��)�Mn���c���	�2�g�,�����hO��&{Ѣ
�!�Cw�a���n%�4���U���i�nTL^�o�A.��.a�˙q�e 9d$w=�I�Ch8)����yX�EMQ���`�R�9�/�Å�yE°F1�3��
,5�V���Z� (y���Y�P������B�`\�̀��}(=�y�c`F)Ӝ�Rr?��F�|P(T�+�)XQ��r�X�J}� �fAHv)�X ��x/���\ɤ�Y0���$��D�B-fE��59��d(J�F�6 21�Z�\	v邍�x���@�p�_�I�X�h'B��,VHZ�Q_�Z%Ȏ�K��sa����3��X�0�[1x� �uQ�zL_�@!��(D0v)�*Z���h�w	/q�c�	U^]Vp�]�	�h�Y�^�9���	��Teː
��	�Z�����Y�4����Y:%b�T�!�1(��>bf��K��h�2�~8�!
�/4����N-�t��K�a�r�Jﰱ@1]� 5!�a�`�I�ֻs��FEw�{7O�R�y&��`�����œh(~�^��_.h�!Y����p_Rq�,^!W��=�Wخ?Q�d���fg=A�Ѽ�>V�N��\jB��/�B�p�N_
WO�?��f��A7���Wl�)n��X���!�\ΫX����J\��[���a*.+��p`Nq)�=�dC���-�l�]����&�CxT]h35���̺)�*V��m�_^0��Y0��k�:��n$�%9^%� �S�@��\Ӯ9̟�I��NC��>hH�����Z�ȿ��9d?1�od��
�PU��.T$�,���]~���h)����w&>Ahnsbj�6�� m�Y���=�9�K�A1ʀ���QRY�-���惞��_+�J��O~׀1��Ql�$�2KT�$*?}ShW`�W��/&�"?̒'YCߘ�-AN���/��	�\@�VAq ��cS;1ǰ�)5K��R�=[F�.v���P�,�v�	x��c���vH�~
q��	G�Ͼ<�d�qp�P��YF�C�-"R�[��u�/^�9�f���M,��-�;�	�7V2�U SCQ5 8�x��@�|�U�!G�y��=O��i�I���/fG���	� �-VP��p�)M���3Yl�Ph eĬZW�y|�}KX��H~bJ���L��Y���9�����kC��t���B�O阾O��:��ր�.6���K�*𳋚�/�a�7&����/\�f��$�W| ��v	B|���xF��<�k�RX���9:�V�&�[x�@�����
����^��PL� %~SK}���,=�z-�����2�����c�ȵ�A���qy	/���~ FZ=�#��.���r����]��[W$΀���g���=Yr^�EQ�n? ��?Uh&�u�jG<bm6@A3�)���ɉ�x%��Aj�z \1Õ��-la���a��N��/�v���+�k���@J#����N��g��V�ع~��>��;7�G�^�	�)��Z�>�O��@�?k�$����|Job���v�	��؀�/K����T���tKW�V5�{Df�u��,Pg,/�ZX!H�0|h�R��DV�" i!hQm/eZ�H�U# 	���.�W���Nd��>A�s<�����P�?��D�ˮ������N|�};�����_������E��|Y'���U�Jy��R���Ceǐ�n�z��[� ��"yd�r�zX���J��H�7G5QJ�T���Lc�%)a{0Ry� [�S��0����g �)�s[���.�	j	�X _�N�:�}]&w�B_Ŏ�-r\,��Q�IQ�5�KI�>�ք�%�8�S|��0:�e���j7HG�B?+�����x�	)�][[�� ��, �Y<�� �/R���j�<k1BX.��i��l9���M{ -Bl�^'�ű�E�Yc-o6	���#k�"�����J$�N�8>/f���cuz��O���a[����LYf�P#V�	� ��A"	.����H�d���W� ��O(D���� !t'�}	#-�ie� ���b�P�l�0zZ�闷�d�Wh�I*���Ry�X��P{|��1��q�	%�v ��!0�ˏI�x��m�YL��MQ���i@h�j\X� �*̣!)���TA�'��z*`�1U�_C�?�eNQ�̘:��~j2�V�	��=Z}*(�������+�����[�	�V� �JAq�&!y���k�|sOI�+Q(1��^��}H�����1���h���	q[����nZ�R�W$���w�[a4���P��[�;ݯ�݈C�2��oԄeT��PXj~ �	kpqBS,<u����+jL�/�2)�� �Na�D(���U^ˁ�����⪄�	\h�X.�Y�Aram�V/oԇY4��Q
�铼P77�z�5;�"����JD�W���W��RQh�H�c�3Q���Wf���=����zB.%.�F��JX�н�°���Eme�����s	�bFZ���51OR��=�"�n���Z%Q����(м�y�%T���:��%�iXeK%�*A����
��K��RAH�ԇ%Y��_VS!V;���O���QPfTX�Sc��p7��j`�a�1�LZ0Q�� 5pL�*x���<>��b�R�%X8C�)�`_�@=�0.�"�9�7CL�����#]�:��Jh�?�&%W~�:of�i��*�����H�J�V��ɦ4T/P�x5��<��m����hT����A�^�ä ��3��]�_me>���ğĭ��􁒮1/B*���Z>O%)�z� ����;!\��	T_�K��X�h�d�I�>��p���$|�VX�QTB��_���>(seU��\�@��,C����ڴ�iI�Ҧ:&�^2�U[�a�}��X(�w����Ē,h'`�N���I��h�):���r ��q�Ԑ�;��&����1�<^U��k�q�a��@�odJ�1
Y�;�V��r��)�_��i��%vJaSx� M]�(K,$	0��2r@&H;�	�`#��d�1���L�~�@0���h[w�z_���X���M���7�\� ��8vd����I�m��6*=���2��h{bM�tĒ5�R�,�9�f�+JX�+���%D� �k�̀��P��T~Qti��=�2S�6%�J�Ż9��@� cT|�e$)��-��x�K��,�XQkڨ�_a��S��z'J�������Y��'Xr}�.�� P� N	�0��"@[1��h�^r2�9�r� 0�x��Y��� r͘M	3�JH�$P��ó��H�'h�����Ud�5]L}�����1c��*+|'q�XfJ�\�%b�`�x��hxJ��g;�\R�YY{t��JKA f��t �ax^��`�?��D��z@l�����P(�X0H�K���[���N����%"W��c��^����9 r��;�p�nIh4��>�qy,��`2�O���������7����"�G�� 
����9��eR��_
�>(,���r�VZ�O��eN%�X��Of���c`��yf	 S�R
t����Ds�����ykxt�7X��c��d�ƍ��X�=Cz8��,(�j�Y�2pX�1�����P"L�Z�|����8�(?ڴ�%��C���0��%XS[g�Y^��p��+܆�6��ǝu I�J� �hX�8�R%�[��y �nZ�E鋲�D�;NVP�7,0��;['��j-[�����h�\{���hM�{)U[-�_*G��T1���K�^0'��%F���$���5t1br?
e�=�[�JJi-�]�Zjȏ�G�?%u�ܽV6a�H�/*��J��#p�U$���b+x���@���ݹ�[.��s���I�YN��ʻ׏���F�Ns,#h�j�
�݆H����*fi'@������w2��%q����g���A`0ep�m��{-a>��X=��^�B�Ag��@�m���2ZNTZ�̯�Z&�b]u1��*²hXm��>'�[�g� =^-|$o�m�xI�d!��`,���V ��^�k��ǟ �kho(]_��mQO��8�$���
v�|�]�E��b7�h[/!�&4v=��OӼ֔.%�`��Ȭ� ��fR��� �IZZ��U�����u=Qx���3B���~�,fXQ����M($�j� � 9)e{���3.�Aw����ĩ&v]������|�&�L�D�w~%���^]�w � � ��{1�Y��$��j/��	1h�z~�d=��[d��R��T /�xeHBv4�8�k���U$�\`��	h,V[3n�B�l�9�&�@� a(��%�D�KY~_�f���>_�H�/��2��hX��^��r� �w'
�1H�r%-�,,���Z���s�3������0_�	%�)t�L����*<��5BO�$�9�PbQE�YA�K+�(Q]XxA��aJ �CX{���*_�/�	ϙ�tS,za�R� P\@��	����z���b�@�Y�2c6��:���Y�9�{-o������?X���DHVFJΉh6�(+$vїF����ޮ �_!�M�?#�	� R���Ҁ�
���|H�� ��/�1	Xh�nt�b�b M�f�I)�X �h�L���c�Q�-���\����`t�	`�CTr��	T_aS�.:Vf�tna�[�wK8�L�t-e�.AH�w��p�µH�nF�	�0Dؔ:@͈r�,�[=0����S	Ks�8(S����J�J6����KM�Yf>�:���?v_V��JM���2i�-$�P�Y�����J�t��	7f�(P�0�;)�3�x�]��g�iL~�%�Y̭�<@4�_u��y!xl��t�R 8f/�?���Í�O6��`"y�F5%jL8���Ӱ�
�C%���1�	G����{ra~Fk� Z���	|Rbά_���D dp2FR��
A�)�ZP���Y/|�j�- �h�/i��&_Y�Z�� �����B�$��B� �gQ�&�S��)!��m��4� ��-|c�"�¨������Z-{َ�zy��_�U�\��M/I<�<�T�h�EU09���$pG{N܀w��,46Z���� gm�v!��`#�5���n(TY�#<%�ؐ�@	���� �#~q�`	�NtP-l߈D%B@4k^(8d��7��x�Ɠ�iFɀv�E 9���	��|~��}��7/V�ݔ*�F)*M��"��ĦX�����U�_����h�ِр�X�|?a�}{)��w_������E�h��l�F` �������<��U��DJ>�{O�i���o���LZ�hI�Y�OBC�����? 75�)�v��'���hD_�j��R�״w�o�}_ ����q�C��젊�r�,�Y�*=��\1�E��5M����C�\�#�=�!�n�8�~t}s�!d���6|��cI�P�8������?V����n��BN��KI<��֧R���%������y��Pc����y��d/`��{!U�&��ry�'f����F�u[f��*ح�,�h��Z
�����2r������ED�v�C�u�z-�R���I)#�*�U�[ ^�9fOK���S价}E'1���X|�h%XWN��X8dZ�%�:�'5@�bኙHp�O��(b�bhU��/P�"A~�7tu/�Y��a	�gj6	���0��3{.����w$Y�	gh�o	�l�",}��RA�D1�R�1u7/"/���y��)T�ZYV��k����o ��V��D$`C�:�AP��G5�g��O���,��h{Q�T��9^�k��>-MFk.pk��Yw.�!�t�0ԤɻP��:szF�
�"ʖ �Rp�hxM�\h�d��qٮ���FF���n�ƀ�o��"Y���]Ѧ@�>m
)��,5�-�V�^ h�5�0�EK��oLz�	��[bi%�dT�,�j��)@a��2i$�H ����?;���s(�m���	)�:�/�jbܠ(�y�<ņ!���G��t:ʈ��
sQi��Y�
	$ѩ'���<� �LRg�[��	�̀��]eEZ�lNF�q0���p.Rh���e/ ������h �� [�B���=�	aJ�I\�v�`[s!��|(���RS@�h0��GP����X��&h`/��*�N)�tX'�����҉���-5�`�b?�"���'���[��D�/�1gWT*�~��e荤ۋP��@u`�6vj�*���[��*Wz�Q���P�� I1����Wawj�f|�� ׊�	�Z5��W�X��(M}���h�c:u�3��lH�%w0 �d���r�L�J{�2R�i�����|����Q����������ׂW�Y�s��xhZ��L�aH�/l��I��W?;��鰤�]�#�Wtč��$�뭄����p)���b;�C�'HO �x�1�^�ߘG�T�=����L�O�""y�a����&_7S\�)�*]!d����5_���yT���!��-�[^���UXv(}�U)�o7~�����/�C9�����F�h�V�@��=��pR�ï��� ���VA��;�hbQ��>�;�ۡ��l�[)��[��hy]�si�r�M�S^�K��!�^	�������P��� ,�A��H �M�	-�E�Nqtz=���ZQ�a�$D X-+85�s�u^�� =� 9���I^فPhD7>���@T1P֤�п�H�9��ˬA� T�'s��`�a@����*WQ�	�6�~���3j�ݗ���X�IG�� �5T�r ��^�VI)�d=������\��%^ 3��-�>�K��©������S� ��	+-1"�XG�	�?��Ҽ����$t��_o1Q,�)1C5�zeJ7R�:h��h��4����R�F�P��%���P�����0'J�z����aj���.HY@��L�%.y�=��pP�A�<Ved��Pݽ쓼a�*�	F���Ɍ��*�n��\!g�Y r���Ha�E��Җ�^K���m�0j^F�0�X�h	]��Ft �{?�.�P1���Ic��V�'q�o�OR�A-,s��煖�����߸��]-�D	e���*i��JVM�Xe �'�6>���Z1D�L�b��`Bu���N/ RhU��VJ���kz4MV��^>>�𖇓,;���I{s�;��[A٤��u@8�`Ud�|GZ黀���)�5�)P�e�K,�9}Q��:Y��A�@˔2�L7v\Uܥ�>�� tG$1�]����F`y�9t�Z�ȑP��l���#.\AF��0�A�+m3�E�m���n�E5,�28>���0��l�����K�]�X�i���';|v�ж�*P��Y� J�+ݵ(,���s��cp�`>� w%�)�3�O��Z-~B�U8'QT������]P����<$r?9�B�X0��ȼ�B�$���(�XȷlY�����d&�A�QHp�
�(q��Z	n����|�h��؞QANe�OYV.6M䀈�'` M��S|zH�y�!��-.1��;� �N2���"*>���f])a���B[ȱ餝�`(�u��^x�����A� �.�vu\�@����0!��&:��Kj��K9�m%W������1��h�I�$��I��sSu���T,���ߡ��$�q$/FF���K�^�W9*�6���|Z�vݚ�X�S���ipҌ^)��z-����3N��K��ZȴG%����|?�6	��!�;i �p�x���q/~ʘ�X*?/R0�;W�����Tղס�h<p,���	ZRшH�$P�ީp��8fQ����G+,�W��X�f�0�M�b\`��h�OR��y d7.^����O�:�~i��:�"�`b�>bw��$\*�	��Q4<	��-VTR��]�5<�8��U�h .���%��@��7_[0#h#�UΑ/�Jׁ URW�:�Ǧ,� (���1eu!�P��0u���I6'����u&�B� K$�G|Gp�h�T�-g~$��Θ�zQ�Ayg�3;�<�_V��@QQ�;)Y�/�-�Eǵ�YVL'�-���^�쾘��`%K e���@�#���I�q�K�3CD��ġ'��Q����A�u%*Ά`�f��h*�(|�*PU��:sS���w�'��68�O��\Up��ͽnҜ^B�_]�g����+/��&'zN`��P��'f��������V���l�7����o#YS���AO<o`pA�{z�=� N�c�Qj��[��V4�)�2���(��`.3;hJ�6]�V�,��yl2C�zK��q��&Xo����q����џ2����B��K�Vd��R�q�A���:��#��T��
�[)���ZC�fXs��O~�9.���:�p���H�ՠ0�X�֚m�L�[^(A�N��*��(�q�;��ᓟ䳶�'Q�b�Qˉ�v�&DS�֣��h%x~��X�Nk�����qm��Ƒ૸�YI�L-�p�u炃�0XCJ�X������ś�\�V�<�^~�����i�bb��h�]9&c���W2�M\W��ۤ~/�p������Qc���+0M����a�:1��~"�9�l8E�~Cy=��/�Wx�w����R�I|�j��L&!(z� 2�����`fh6s$�3>�F���||x\oWT�C)��^V`�"_��`0�&1�#�~*�ni�E��b��\*�v�(J�UT����C��̱<7J�VX�$����|Lq轗�#'Y�uާ-�<��%q��hsK_��C�	��#��Mhx[k��\$-u|^�²���oȔ(E^$-�g�w>	l��"u:Ȳ�P�q9;]~ѧb�����.�2	�
FA1�q��]� �&"�n�bB��D��	��'A�XW��Ub�b �^��!'GL� U|�Ω�Z�@(��e��������5�pi�y@Q8F� .�h~P��Z�����H��f�aJ`��$N���<�@�׈<`������ ����%��X �`�^�eM|#,�	�a���\�+��Jвx��q�5w/�@��I���K�J�����D�=�|?�raක�k��{������1l��n������Y��?���^{A��G��`�d1��@<�/^fH�R�0�0'��@.�(�A	%��0f��`%qt� �t'q�bf��V��zk٘/BM��3OmK#�����*�5L[O��J�A��Yj����k�A�J�i��o���^T\�h�y��j�	7 A�1@��2'�笗eP����T<���#���-�<l�SIEPT��Ĭ(�Ү,O@��j��+�]h�����/�*��e�:m��)�E��� �z=H&:~	bMC��LP)��T�Q��ÿ�
h
�ǯ��&�+j=�����]ض��x2qa���)���~��>�3j�XԀ����b	�����h��a10�:ȠEY(*��/y��/ب�`�.��` �{'�>�Q�9�x��
{�^yrp�1aը~SĽ)�\O8���>V�61X\��>�3��Qh�%\�b��$H$-� �Zh�^�#Ss �쫵�	� 0���at�F�X^�A���`�AF�P�^�SR����+{�v��:�G�`���4�"([,��to)`w��9��]Xl� ��Q^�;K�� �52o�@ V6�3���p���U_<����bx�ϧu`��W��L���)�MzZ8I!��|��>�N}�r�fw�Q�w \h�b��*��QS,��}���X��P1P�c��qhU2���EV���z?�����/^��;.mF�ϻ�}�-�L�-�y+H��vO����]q�9R�t��u�L�E��ܬP��%B�����eo'�\�oUI�-HG���ĕ��[)�:�˭p%� �V:��-9:����Q~9e!ɾ�T]�+�E	օ)��Z�4���v�� ɞ?8�C��j�:Y�2���UrȄ���~�0.7���Z�)<*<CfH!��uv��'B�*�����9RXJpW�d�L2�@$���:�	�Z@�l�Y=�q�7moi�TY���Q�����{ �C�A&���;}�u��k^�8���>�G�����yP1g_��-+�Gn#
�2�j������x�_�ʮbBT^��x,t��=>?�S1 �eIA��P�?�����K1�Y�}�NE�)a`�\�A�&���b�t�fW �]�5�_���9h_0s��OA%���-J�@�P��qg���W-����_�Z*$ǌshyp���eۯ)�~ �j�e��`�Z�@��i���R�YP��eK��s����t�h�����V�������;��d��q`f}�,+�K�t�iB�� �/�&-B|�+>B�iB�hFTebd^�t;(YR���Z�&����q�E;�WH8t_��+��`	�g��l�]�j/��`|h�r��˄�T���9���(� ǁ�~�\L��{Hx/"���I�(����0�%h�K@�R�Q�c /569�#8���w"�@(u��%�Ѱ�}&��J�J��l� ���:����Z�� -9siO��ї贺�@X_O�F1y-nB��
f��eo(��.sT�f�p�\�x�2iL�7���iI�	B�VkHr��N�H����{�"��&�3�T��!��W_����el�'Z��:���������29�>��r^U�[hcH3_�����j0l�'E�EX_RIV���-�����t)R��%/N�x5�䩸���*���*���( 2�N,���[A$�A��a�,���"[�'Y���w/OOӉ݅�3�)�>�$\a���5q]N�B�0�V�.��H	("�`YzwD>|�a�$I|� M��Y��^��J]+�\P"��޼[P�D<���-S���!U��|-�Ҫ ��h�0��.7� ��.��	�NW��)HRVh�(7i���I|bvDݜ�%h�T�;�Q)	t`��Z],<A�.�:�C���7 S�#<*�>�:ۦ��9�G��p�Q"�J���� d	�t� �o%s4�)6�|�U��a�/��H�$Ɖ�J�A��\��]5��,a�.g&R#ը%R�'ז�дb�� ���W٭(�O�hP�de��E4[�� ��^�ah�S�"5k��������^[�?�bCw/x,��]C�K朄yZ���2�0�V�#��[��k$�	�媻�[{m+W*-�d`����c�	p?��^�5�H�Kd֝dhݐ�-�Z�5��$(VA����;-��3�
��0?�[�������J����?�Q^�Z��	�߸thZv�Ĕ�[f�L�hDZ� `NP��oQ��&1�Xh�
f��h����`�����A�)�,����,T�	�ߔ�������n��b{-ƉY5�+�h�'�������z˸]f�/�KQB��J��Bzs}l#�Pc�! 
�'I�:1���w/���%� o�V�)[>� L�m��x*z�Ha�W�V�9Z~x|�T�㹙ॄe��{���FO���(Zh3 ��������m���}.YQb���\�P|@�)w�KcM���r�Wl��*$kp:c��-
�;��M4�B���~mt�^p�3�c�4��b�@7[�IPhBH\9�W^t\�`J�Z�Avi�q�*�ٚ�E�1��r��j5w̌�����Q;�Y��4/6�5	�u��8���A��l-HrJ"�o��Ln��@�2X���O)�u�1���h3Jp�2%��B�Ͱw}ϼ�Il+[�u�5np�dq]� P�Z�PJ�2+�.��ZfX�v�z� R��ï�q��;!�K��-T�O�	Qfw�:l��1��P�*^���j<�F��s�Y<7���[-L.�&%�I�23]2乼(l�'RۄEZ�U>2��V}b/֢i��|*�'���#�+o��A�3Hcz�"¸l����i� �|	b�w0u%��Љ�_(Y� �Z%8(�%���\Ye[�o�N�Mꆘ��|�)X��K���(ȫ��,U����H� �p)�}����Aj/l���娑�{>lWp��2�.��cPK�w�/ �}��)��JZԒeY�<Ar���*�J��-�^�2�%[X�w����c����*���s]ˢ���w��ߙ^)�a���`G�,�1L:��ä����
zO�d���";�ⓤ�~^�1$<;�NW��{5���8��  j'(�0�su��X��i�N\f�����ݔ7������p)���P��X\KSQ����F�O�����W`Gh9a�	�o�� OQ�s%txr��(��'���<�`>�}�6	�Y�xC�sah���k�a�b	�"�&O����fWR� }(fP��T�9Ѓ�2�F^|���P���<5
X��RҒ�_�]v(��mO��<O�ǖ�\���@h�J����f�����~!����ֻ?���R��S�SN���b9��$�ZTch|c�EH�j�l)[J�L
Ÿ5�Ղ/.Ƅ��8�k-�3 )q��O�)\t0�U+`YX��G�{ra���vHT�Ac�F�TJ����9�΃�ĂG�)�*KǨ���m��u0h%�2����Zl��"q�+�Z�\UU/���� K�\	�gj��h�\j3����g?��XZ�PA�!A�*f.�:���wTZ�K������(���l���HЀ��Q<�`�Jr��^��#Akej(�-}/D���8R�{^���C
[
�����[�h`�����4������S���k4�R��B���4K!QhfC �'ř�K�V'܇p��-��Y���*(�D��N�VH��:@��S�}�N= Z-�/(�V1B���>���#-�S	F��'-��@�1)�q��Bn�J� �oV
��y_;*�v}~�E������zsV]'���P��ב���Vx;HUq*�ӑ*�� �ohs��P �Y�/��G-�7b��px��v�l��	B�w��B%]�'p����^ar1y.��
�V�Hj�����Z��p�h-\�.�NsR��Sn��?���th(����LxL`�IA<v���ad�3|�}^#���P�-�r��za�f(���O������y�-�#��d4s�ɮx���LU d�62/�:*��,<��9P�=��z��A��/C&�����E�*�h���%ӹ���\������Z�Z�&�À�!P ѻ��0�-Z���?"�(��Fs����A�db����@fT�Z֦xN���J�R��E��T��Y@�[޾8'�۰�`���x?#�0�1�½앗8����"7H.P�P��?3Q����`�t��JV�օ1���3��*�����l�ƧcD��.�Θ�>�uz��OG*����/%T�@�=,:��	|�R]&�Y�H��,�m�0��PuRJ���@y\�z�K4����^I��v����4r_��LT��� SWh�r�_�ϼ.,��s�>LR"sL[�O��K�V����;�pN��J�Oc-�n���i
�J�Ӂ��6dCp�j�w�k_�む�jJQs_��=s���0W:�u��-�b�}��%�3�Q �׫��!u�-�Id|������P�>!��X>���A��_Ah��Q�g�����-0��餹�z�o'QT�����] �ـ��0����];-ӥa!p���h?I�|$U4���=�:K����A��He�4?�:QZz��%��K[lJ��4��^A�_!~�� Y	���Y��sCoN�B_�3'���/�^���/x#�U��%��y.9Q���ץ��j�a����(<�,��K@큁���;!��[�����)�av��0.�~��*�ݎ��D�TW��D�pьS)���>�ֈjs. [�O�Hh5�Y�/L�IT�����qP�����n�v���oՙI�Z����@ؾW�a�!����QL��(AE1v��T.0���]*�t��.��ź��+�#!�	�TZ'T���a?��d5(�Z���J�
h^�b�%��P�,0�F&(ح�v�B��H�50�{w��
<F5��"�Ѣ�t�¥��)�ъ����zg��o��Ӕ�&Z@-a>r ��h\`V�/��@���7\���G�:,$[��A�.�۲LFt�p�k7�G���>�V�	�/O�4d�7T�\@u'Y���YGA�nXh�KA���.��Y�jc+w� hx�&uU(|,X<��xx��^> ���m7T�8��O5@Y�,�   ~4H6	�g[5�nX�A��_��h9*-6T-�ZY�/	�ZPn&�F���,�O(�)���p��L.���CX��'��P�<�ȑ�����{!�<�=�,0�N�.��	�;���/ ��l?�g��#'�c�$u	G�vZ�"��`���#|Lz�g��]ਖ9����J	l~��(��
�m���2��o,�K��誈�g���p�#H��^�JK�)Ď�ҽ��ж�� �?�w��U~(�7�<ND�{t[��w�	���֘Z!���:�'h/os� ���0�{���ZNd�rto���"�O��cS6��韎UDzh�ri_�h!;� ���.d����6/*���Ps*!���*�P� =4EV�� ���"� �{P?wYsL !$F�x��&�t J�_N�q<�@�W௄��k�](ꀂ-�@d鲴  ������r�~M��H&�����1�)-0gbH��_UW���'���&5������ݞ(E�%Q�� %�7�5�3u���S�ۿ	��b�� ���^��:'��GǴ��>�_,��E���p�V/F��]�-�
ړ-���2A� Ɗ[[3~QѺcf�_���-���(�Ů8�l@qZ%���
J���p�b)�'@���葦�:�MX�v�ް[	�}��W��[��9��5|�`T�RS�v�PÕx�,%`̅h��rH�֭�I��BV#�?��#U�E���)�y��d��0*!w�Ұ/�
���xr�r��%B]4��	�C�4ߍ�?���Z:�l�Q��� �m2�*w,T����]"V�A�%!?`6�-_�@F
�&��jW����ۉ���;��&yx�T�X0��Չ��e�Ď"1W\H-�+r��_&-���?�0�L�iwm(�P	�yL�~��@(�ـ)�sZ{���3� F?�x@Z��Җ����c+`�e�0��M�#��J�Db׋- 	�haF����e� ���GRt�!AA��BifV�d�޳pH�� @%=w�5# PZ����1U�z0�C�q~.�}�xE�q^yh"%|Nħ�	S�1�/�\��S��\�X���h�=�NJ�$�)�	��[�y��8X՘���'rp�*Uq�@��5Yqh1��u��T���Oq�:��y
��Z��p&1c�n��<$J��P@�ZM;�`	X[@Հ�51	�i�ٕba_ �!U\`y	�{?C���8!/��[�-w ��~j|*8���o��_�&�
]�J��>�z��0+W���V�rΠ��I�$����(�A`AL�(V� �@
�T�kIՈ�$�4 Ph.}�X���ca�P�.��2�X���U�H� ��XY'����`�]ӧ�{a��h�v&����0�B������@{!*�9G�/�+l�Ų����R������9��hNs8ӯEC1h����eF�)�!־q�K�A�E1w.���.�a�u<`�Y}�'̉��.h��2�X}1��H��N���=vU�q�R�ȇ�1�(�ݽqC+L�ĩ0�CЖ�-m�38;�K��+��)Oe1ϑ���p��%_��z�������v����s����TnNߣ�A	��Zs��Hh�YʻlKW�lJ��2��5�W���j¬�[b��}�[�|zK�(�&NR�-4웞9�h�g�4[���UN-����o��DP ��� �����B�o�)$?+�;�ި9fP�IJ���-���h-�7ٖ������e(�r���h�w�k���a��҉1%1.�[�E<�{	�S,Y�'$tO���I������	>2,i��S��$P�h��& g��ql3���[= 0��!0�t��9'�ˀB��'�1�pBH<|��@;k��*�K��ѓ�w����S��Eny�BϘ՞ҼoIP�/餆�OF~U0�y��cy)�� �}.]��E-�߿�p:����4	�Ar@M��fNX����[p�K88�vk�H%�'�0</Qj	�}ea��*�Y'!�$��d�4S���X�	�3�I�%1���Uh3��K\]��:E���D���_͈����W�$� �U(�f}YZ��@X#��x	�EN���6�����g-AS �;m`W�6�'v�ď�d���JN�)�.S���:	]Pt�$(�~
O \��h&?n\��R����`�X���#0].$r�^Y r��,�(莟̿W�6:)�Zp[B�c�T��P��J��Y��]	��^8�d�Yt8t.���F��K�� �n��W8XF^�{�D�>�9SK��U]���3n�1��X&lQ^���B8�m�bTુ��)��T�ߥ����| Mf���i�)ֳ?-�'����m�nfp0X�_�E�3"h�`��@��2x!࿋x�H1_&Z�z��d�r���yIn���� ���ā��_Y`����px�n�Gj��TQ�Zb(t�~�;��i#w�<P���T�%}WQ��q ��9-�.��ѓ�_c!�K

�3�%�45�/����:��'Į���<7��K�!O�/���d@��#�,���������~S�</J��9��*�ߢ�V���R��$�¥��@�x�P�;$]���d��V�Y#h�q(H Zl_��fz.K{��I	����=$/���uJ�9�	� c���
���L�
���p}�u�pZ�Y,��hHT/0i��M�)+8��E��P�"�+��V�C$�x�;O촉�yB'^ڬ�Z ��/(*��L	=81��(p�*�@��r�z:���:��NMt����$2�X��.z�0��=L)h�R4�ܾ�M��:30p����
1
�R<H�	h�,j� `��N��� B�%���~�R^ݲ��Д\�@Ä^'A{�7h�6S\������?D�)����LG�~J*�kEHjʈH�}>�?���fZx���4ԭs�NB�5�4��	h6}U�H_����/����b� �������d.QW_�((�?����7k�.�Ϙ��}�I�H=&�	|V�m��2�*>%\!��ƿAv�>OBL�^�&j�X�q%D�LU]�\U�TL�Z��P��8�d����E�e'�#QͶAw�I�g0d,hM[3��[�q �N��U DOF�yK�� ��n�A��p!-�[:,��{J�0���K
�����_�W�i(�xSv�w���ן]{, o��-���%���H1����O�H�nS91�5��̴���N���,#���:��.�;)<��B�]wţ���/���n$��V}˨hso��PiZ,�H�u�Aa2����j��a�X|Jp ��QT-�� i��Y1�_&�q�����s�6~ ��R� pI��=�~Z����o*jn�J��ƣ�H�^�� �0�\u>vHQJp|�PYc�A�z�D�Je�?m^L��0S�'%�I`3MT\e�C�2^�y�ZQ�<��ǔ*d����/�Z��,�e5�.Y}��Ȝ8��]�5� �vw�N���d��X��`�?D3�Q~�v����X7OZF���a�����y�&g�iÂ��Z��[T�����	ԝ`���a���~�B-��L�`>�n *�.���i_)�$���+�y8�rL=8�7ӠSZ(��r~
hXݼ���(E�4K���
`c ��(w��t��/�̱.����!�J�yM��}�w�Bo��J ��}AEHM]��:���1��t%a)�� ��@yX��Q��g��Y6K嫌����x2-8�٢D���!�sV���`t�T-��c��^�_�)}j8�0'n.h�o���]��/�bh�f���X7R�&S��q�OA���>��P�uRQ9���Y��F{��&�'�;�e��p�'��� }\�e:�H��CG���BV�d�11�(x@��%N�U5��2���{y�D�D�ޔ��+N�/$"S8���	�����i�X���0�[߂�	��C��S�����P�L6(o��[}��SH���2K�Py_�O��$V��E�*$�F�UJ��B�����rr`)����F(�Xh�qFB[���%�k�Z�K�2.5�c��w8����UPVX�J<{vI���E�߄�[�q��hDQ��q/@0��L�B@^�s�	�XR�_!�j	����(���*x���v��_��+�KH�i&qaI<�oȘ�f j4s��1���c{�w�z2˫��Im�`7�?����7��8jV�ld$-	�*�@�B�W-I��P��#�X�0���~�/�d[0���l�Z�6�l�-�%C��Po[��~D������^o��RA��r+��%w��U���(k4���82)ڻ��a�`���+�}�n�^ZT)�@��YZu�#�z����4�J�Z`B�Mʹ�8�IJj<D�TX��M�H��&�)�闁ih��pHjˀ���R�N`��	/0�	+\�K��B�p�)2������� ����H#�_�@L��Qه+�a�e�ڃ�~���2'?=�a.�|=v��!ٽ%��� M�E�R�R�1_YSpXb�S轷\��3s����T:�e���y��]089^��Z��O!�� �r�.1�(������Ïh���@���Z�k��6���@�^�6QVz�:�	�7/3~���{[�w"$�/�kE���p����-	5�hz�F��etO� �ՠj��=�8	_���XV��a�A�s�j�)��%U`ýcdb�h�AL�!=��e��g*�����%F�! OV�2h�Rm+KZB��#�H�c���YKy�/�d ��&���������t*��#F�m�ϱeW~�l5������l�H)���a΢j��ҵ$91]�[SE���_�R�,��O���r@��fy_����Gk�qy'��r�N]���m_r�	�:	�W�k�o?��y$HPZ�^�/,ɚE���w01}m�<�9�:-� �UN.�dk�.;����Z��������4��0��;�D��O�Uz��[g0>��.:.�Q|l�A=(��	�!��Xhr�*���4v�k�9s�͒y/t��U݋�tҀų�|71P����	�t�3���@�>tY��A3�ŉ�[�VI>�ih-�1џ��_]��,*�<���Iy���8� #j�պ�?@��X�����0�,y��t��y�>
Z'V��S|�,�����v쵲_.��F���m~K} 
�˂�䘥�j���}i�'�Q��U���=f}�tv�x�B����s ��~/L���pK�ZkeV�^閞�;[-�.��]�*R哥���!�
/�	�b�}�&%��S��>sդ���OWh�7NJ_!��T S�?zs�е�hR�y-�	��|����ZhUMx#��d�"��h��n&O_�V!�_�u�X	�7�pc�aW��Ԁ�5>�p�Nޅ"�)�.�1X<74��H)zO6�[���1���I�4�(ؕu�ʅA��>�Y��z���!��)�y� i]p~�,@RHt%o--(��:�7R�	hj��YA�UO,|~E_t�W+$��|��A� d:%}x�02����XE"^��KG��-���1�͜�����=�d�����F)�ﴠXT�ȯ@�����	{��:$�� (���0v� �,�g�y_KS�[>"����d�PX�"2K/!D�`C���i'P�N�Kh1�(�M�]�>W֕:UU͞	����]����r��Xߏ4u%�hm����Յ�"�dJ��	X�gJM0�y)�
Zh@K"��pXP	�|��)9�k]-���`+V�h�{P@���}��:��� n�8~�f��p?0{G2��F�	q� �=9J��DCi�f�-��^���l]�S@�X ]�x�5�Ð�JQ�)O�4����-�-̇�Sey����4�8��*+���B
6i�U�H.�[S��1�	so#��EPj�.������X_/*V��N�r�"X�I��	�B"�_��`��p��@?5���`F��4���ũ1;�xHi����� ���{�1ϵe���~���5re�}���c�8>c�h��i\:9��$���[Z1�U��R��� �����:^=b�B�2Y1��ҮI	)�:�2��GzfyZRn�pk)x��������.b@;A�w�u��FT�u�N�u ��Z�?M靠S]�>�j�@��_�
O���}=��-E��,�������}�f��\��x���a5Xh������N��Ӑ�(�,��޽�'cEu�R��[�]�L� �<N>Q� bC�M1�Y!��������Ah�z�:�S}_�\�$z��_�-��,�< �MPv��	(j�f֊'r�c�
�_/Dy.�*}m�>���\%�CH���DO�5g8�W�;��P��xqc��H�<�������|��M��K:2��d���P?Z@"�.�=@����W3:�PP����] I�O\
�����-;o�Jz���J�
�6��Ƨ��-#�MPH�x��A�n�΂�Π�h~0�2Z�kY����?�q�E��W�u<$ci-tB�/��V�T� �ttP�J��A1�:��9mjF�]�oZ�����T?��	��$Z���h���i	{�y���K�\�7�A;D\��(Nc�>�1��/��ց�"&�%����XU�΀Ah�,��V�R� �[��X��~9}$G� 9�����K��|��[6[H �ǆ*�q��z�,;p@��1�3���$�+W��w�1q:�k�;,/��� �:(�V�@
)���C�`]��rB@W�����K�T>�`t�����{�j��1�Yblq`�g7!���x� @��03	L*g[���N)�:ع&@��9����F�̴�T�RR��v_��6�������[�чh��Y(�"�w���1� �5H*�I1�1,�h�t�A��(�����$��L�	�Ї	�'�ļ�pf���5�JZ+4���y{�I��V��^_턺�c�yH�rA2�׫aV�}n��mtU�#��t-8bE���t�W��@�K�=���w�v�u�yH-h��W�)��-�P_L)@f�K�[�n%TLpg�aSd���LD�<_����r��nym��f+���X���	Ԩ�T��ٿًX��b�K�9?���ڶ	�EHK��:M5)��@X�w�����R��>�qqdգ�|��Ɓ�d�KR�l�0�J�j-�1��Z��i�ll*)���D� �%|�U�v�5a�Zjs�<��O!{�d�Ք7���0��[�h>�C�c�?Zû�/0�w$��h���^
T��L�(��%�-�N�f|\'��"�)_&;��,�� ������0�e���L��d�xt,�l��ݓ�pT��(���h�KсPQ�c���"i8	��]˩A�{(�Q��^H2��9L�3_�w��������g�> ��)����ŕ1�s����,&�|�N�߫]��eƲ	�RL	�%ٞK"d_O���)�%z�-$��!9�Oۺ�=���fqa<Z����R	Ҭ�*���1�2�T�(fh�PNՊ�|'�sS�h/e�{����6"�h������x�/Y�,��HI+!0�d��N�KvWԬ&�^�/Y\-�.��~[�W�1��{�CVp�]Z%9*"��Yk���|9�" ���@JH|�m0�cX�������L ����R�Ѐ�H���-"��sx
=ڬ�=�F1�>��>m�3�8
y9�.s�`$��.�q��P�&w��c�!��[9)h03_0��I;PT(��Ok�wX�ZH@�ID�L�P޺��ܫ��@�lY�X���^9��[��1�?����pA��i@l/�|/��l�DDY��t�D;9�Php@�/���C$
[�i�F�r�"���h��Pk��
�r�7L-;MP>�А2 T��F%y���@��y52߮K�I��0<�6�j�?B�����.�H��џN��сBE)�����''V4Z�U�Q�!-]b�r�����Id.=���� 1�XS�q�:��Pg�Qe����X�B$4�VB�3w��e�S3�ʸ �XF�_����h�N'���b�{��Iň O��Yah`rs30�2�fR������B�;RW�H�,�'�!�Z+��%���h��� /��$�W��p�Khժ�4����]�À��,�u<5꽴
	���!1A��*�4�<Ε�F,n��������YECim�9�[ؿK�GR�Lv�bC2�>n���S{�k�W����H��y�3�CI5(3U�H�Z��u)$���h;
���F\�'0g�@=�5�}v��	Uғ����S׎���0��2�@?���|�9�O&��.Q��-�.m���h1W��v?V�Oj��[;�?V���gȌ�Z��Pyx'���C�C%$aAߘu4n�r!�,6�KUd`s��܂��iPQ�*��		OUl/1���v:�|L�.D�\ dJ�O�a$w}�HA�%�>w��~���I�_�'s�8-�Bb��F\�m��@1�S��}-�*��<�kN�-��r>�P�JY�*�U � ��&hw��ฅvj1�^���u)��	�e�g ��4�(�J�����q+P�AA*�Op�)�j�}'T���Ҁ��<��hx���m�.�2�z#M]RO�gV��u��[)�8qn!h+,�h%�}�u����΀��S�E��I��L���-�bV��!�H��	��~�T��nBӿfw�!4�,�a�+�WQ�p�=k����}Ph�V �b'
0�u�t�̱�S���������I���W �~�z	�=t���F�<`�H	jx����H��LgW��_Qr���BhTi i�љ ����U�y�4��l.7�0�ŻTB��)����;_X.�X� �k)��KqTbkuqm�}a�����^�zN΄K��!	b8 �C`U��J�i��o&�L���n�8��P�f
�v�Bz����pf��)�򬗏=���4��ž�h#��T�[���q�*@+�>�9D�?	�Tu(5Z]��n2�X��Be_��(���W��0'�z� � S�v�"����wl;�rK�P����X_�VYXހ)���؁�W\4�9��=MLVdZ����l��İ�*��J��!��Tl�ۿ�>^�(,PhR	�F�U���[=�����ᣴc�Dՠ�hQ�Y:Ws��3ĥv��xNTV�6!#��-���*�������|�_]��-��p ��+hBd�["����{SK���'��������h�_J� ��r�@�0	��>���z�[6рKT�ǺWK�KF�vZ�h�����gP��f3Z>0,�&eD�_O�?;�>q�r@˿�'a��&526K�k�נ`wA`~��Pk��y�	a�YsB�� P���8%�F/�8�/f�1]Cuh8p�������*��c�i���wsM�(0�,���i���>i��R�z��)�/b��
!��-b7|�of���͔X�EB�u@�,����v��q	[��ʉ����	��&�(���!�8�H�TG��mWY�ZX�tbh�O>4���+0v �Zm'��޼��Љ���IS��{�!�f7�4��t����U�߄�/� �������z���E�'O[H	s�2��!�؄0�'*Hm�D�?���'7)n弓�t�!�!���E5^����(DuY�I�5$�{pn�_X��ǟÀP���Y��&@*h^�oOI���������FO��_Fk/�W% gf�����H�,p��7�CP,-�Y�O����]/'�L٘�`�P��M�LGO���8UWh+tr�0��k)%LoV(鯕����l���R�?u.
v�N$tB*����QW012�*�6h�l�j��kWaqFi�m�\��v)
	XR��#��b��M8�N좰(�,_��C��C�r?�J� Ѽ:�@���ϻ-=�����+���U:��.��Zaxln7ɒ�THR�pW0�8$=��X�cQfA
Z� %R$�"D�O�5���V�-��)�
?�ڬ�	��ջ��-e�%�h]C�� �c.7,�a�1��*��ֳXFWZ��*�;�*��,{R-e��\�WZP�\�<��5jG���{��r�Nؐ�VYZ ��6haw�/��<4�-x��]'T�q�+ѭ�'�VG�!�o0�s/��D��� �S�x@-	��0(�_�	�gkߓ��q|����6:�_�V�7���erK!B+)�!,|��^���.mHQ�p\T�'�s�a�?j�8����qx�`���N$hX��5׌�)a�q�%��h��<'T�@+s=b���l�{����wu�pt��@��!��Z��	��y30�B�p�{���R����s{��?K�q��젖�T1�0Y�[N%+��w���P���DP7�����R�����	|2 �.�!-�,��BGǜvl\��O04������V�R>^S-p��`]4q.�с-��)1��ݳo�Ip6�fY��!�
>��M� ��W�r�N8�s���r
�چ-�o~5�d��+-fz�.�[B��]E
q�/��^<3-C@f�[/�A�Go�����y[��+X�0�<:L� �lG�C-	krNO�/8��c�G����2,Y�����w�ʏ ��+�rfy"w�^ $���a�%U��h"����������h-fT�a�t��g IN��-���r�]�������J/ ��-.iFQ�V���|p:�[Lh�MZJ�@I�_|0��,_��>:�iUg�\�h}]��B� ��!j^��x���[&��_0	FvZ�	2y� �sزɘ9(��0�r��K��o�bC;��kAߜ��� GP��sBo�Ws�,�K��§��������h�>�N=|M�v0���0��aa�(�����Ed&2��~��W�����0�i�/qhC,鈢 �bfS['�-����K��_���ΉIZ[�`��8V���)�[���-�`�KB_^��s�O�:�Ʋ/�����Ղ4�*��"�l~hIZ4���i��ԑ��!<�[���&�nDs��_��1J֒����6@�h%/d�wl�����i��b�U>d�CV��=f/��FP� �IY���$��ց�Eg�}{�p>AK+�ث���y��[S�O��´�M�	�*���#�P�H��bc,�I�PU�o.��B	�`�K�`{����/�����X���$�>�C=�Z��*�����D�`���[T��,[�)gʵ_������~�21�\��h9*�����ěm	Y���t��-�Бh���D��1�_���M]�HR �Pj�xi��l���z.�m�{�,������h�8M�l��t�R�Q#�`iX."� �n4O��W0M��Q�g=A�Lj��P�� ���P��#�	<�VN�'��z�J��[=�� O���K �(_Y6B�"���ђ������0�S ���-{�~��`�P��N	�?���׻Z{2�l�G��}�)E��K�a��h�w��Qh.3C£�]h�e+�����K!��l5��͒�@L�.�lR�!?�p�VUhd�{2`G���R���]@�2�q��V�N�ƥ�W��H��e,��,�\�C��2`�_��Bz�h�ˠY��t�-�#h� �%J���5N���w����E��qt��q*�,�Da@��`%��3/ο���)�h2D�~��tO&�/Oio���l�i7W*�Z����;¥+_`�Cv<��4�q��V?��A�<f=�N]�+��|į���*����wS쏺6'g�����)s�Bzf�z�TT����2&a�Z+���.!�P6Q�x�kd�q��tL�F��͋
 X9MQ��gJ.�e@���G�!�*aL4S��@�9���&�����,��G��v`��6<-��L8�J�1���x�]�Ӭ+�[���Z��E@M���:� O�A	Rh1�C7L*�b�գ�F���%��"t����0h�VM�-����Ŷ���w��F(�$XQ{���x'WaHR�y�����V{'�V`qN�t�_��%]WURO���)`��[$)�*�S��O��弥�}27g�7���w.�&� ��r����YVl@��/q?�9��6���	��)V���=S��.�� ���	- ��AqT&z*LZzJ%`3�$@*����W�|�M�%^��o���h�#��
c��`>锕�J�xeT��Sh�fnZ,c�V�>`�
�:��+�,ŧb	�"O6�m�:D?lo����	���Ae�Az�h�-��n��' ��%k���hX��F�=�7���C������
	���(u	��Lv�o	_��R��sM@]���_L+вʄ402'?.L}l���Dh�&	�G*�fQ	D]��'H��E���0h�e�Zp�� K��*�@CSwT �-���[B�����ÍQvF?|ar' ���y}950��	��ʉջ�a~x{����ՠH_O��'*@��T�R][e꽜�e��.{h5����mo��%2�3�)��#���غpp����Sy�~0��?�
�HL�>մ�Y�q%�+�|��C
1m��+���Y\U�du����&-:�ŰS�P	H:	Pz��YA�Z1!�5�����"t�h�/m�1�n�^ `_qLN��q$�f���'ne�����Y-�t��A�k����~d�}��PB :0��پ? ]�S�K�+?�=�[�C�lS'�"�j�#�ɧ�<]V�!d_��4��Ni���Dj\/��|��v+GT�F¤���]ѥ?�fBa�RT����<������1	�͔]^�
)޶�@��J�=�%����N����Mq�ΆB���(!�YY'���XP�D�H�j���#l�h�_̯)g�I�r�mVI@H*Y��P�X=SU_��1��݀��}�>&��ʂ�Cs/�`�$���Y-�(�* �N\,X+ �Q-*�?��T$����������6��ޘ�R@��g<)�r�]cc�q.��	2���b�' =X�Ϻ�Y*��i�@r�F %:5wE4�<� =r�mG}/�
�o	^D܄{<�}`�	�KX� W�r�_Ȳ�`"_��2�7�����s���#��ݒ�w@S���@�
5��b�pOw��a-�C����ɜajf/����C�ؕ'��<�(���h1:,F���Y�,�[���-�h~	�W�{	���姈S�B�� �2�c��Ҁ5�"~v�})EB�%h��\B\���c@�0{�K��;F��I�=��{�[y���j���a�˩ �aH/�s، �=H]�&TAP�N�p��2��&�)�5@Y�S�P�'�/�~7bh_϶�'_��R8�OJ�R@Yh�� Li����)K��dN��u�N}��siq�vx,|�� (2K���E-�a�\Z1�{���l�H$ �B^)�Z��� �O�\x�@� �zD�	����^���ɤ�}G����U�JĄ��~]�yQA�V���u���h*l�`�"$�P*/s߽}�v݊�u����p�_A��DXF4��{�J���T[V�4}�����䠁 ��-h�~�o�+��G�h�q�<`� *-
)|��@cT�����hEوߴ4��{�\1��A�T�%W��X��l[Wu�)D휻�ރ�h��|�_:�̾�g.)�蓱Ƨ �>SE��X �mt1K?�F`�:2����-w$�92%b`�g#�%�ŏ'G>��gX����g�fń��U
O=���Y�q1�k�w�zԂ�t�MP~�МA�n��cJ=��Jd��u�" �����,UW��Sb��I�� vS�'����du��T�nOh�e_��t�y����׆!��(�-A�"F}9��`9�Or��@�H>oKt��_�"�Zז )��I�2�z�O�%e�	�5\&��Qŵ�=O�\53�x%L���hE�8����~�i�.����_xu%W����Q'ˀ�{�b����q	�-�2h�ڹ$������#Ubc+�VkD*wr��J�w�U��W�lO��؅�������mw]��'((`<Z�RƝ��"J�AIT]�1T�ѿ?��X�Q�M�q�o��*�S�q��$�2!V��b	�!6d���D��2gyy�r�J)N<�ᇜf��h2�ߎ1�R4�ħT�f��EUU�K���2oqF�e��h<Z�(�:X�O�}���a�(U0J���]��~��tb�	}���7�`sH&��1�Q�z�v h�R�e�6�r�-��P��7xg=�EKp	 6�����hHg����%�?�SQ��[�@8Ϥ�K�p�+��K�TO���A��<�"/�]Ao�O�L�D1��	�[��$%���s1l��~崃�KS��������l��SX��ų����V� �\Z���}�wg�!��Z�ģ��H\�(�I�m^�&��TJ%��u[w�$���UJ��~B�}8�]~���L�wZ��]��@�p�ö��aKð {8h�1J�SW*�.�a�	��}F�{T,�Q"��Ql%"2��)�HXttX��h�78��ds�t���I`x��_F��� ��g�SO��o�Jl6��Z�(�@>ZWh�(F؟ZY����lH�	)r���h�"%Y��p�	]M����)b 6.ɪWZp�LGa�1l�Dבg���ʄ�L%:<ވɂc��t�Z�F/ϩ��a�Qpli��0뜠�h�_�[�a�8`NO�����j=GQ��@T��4���,~�	���P����]�Ѻ,���)���(��n�{`ށ��j'�,��h��`�+ɷp�/7,�L9b�bP����Y�7Ո�	ZQ]<w�������.�Ba`�_p���+;xsi��!�_�"���߄C��6���$����-�j��,G%}�
���$�P��V�tYR~�iBMH8n�(.-�ǠYu�/�p�NO�YI���K��i�Gȯ̈��\��h�JY�x�J��J��/^7�ۤ�K�
8��͠�ǎX�����vi��UG��Pf��|�)^�0 �g����,AT?��@�K�O�!��*�� Ph"� X��%R4G�i�^�^���	�6�Ҳ鯅[�6��OLl�Y�B�/���&��dL����
h�f��Ȳ�K��,� �f�#q��\�mv����$�?�6ob��%�������>�"�F2KoѨ�Y�	x����A�Qkʽ���]���ʀhSO5��wA�:��ho�t�c�?�\�T�9�ep)*��Z�C;��^X�*�%�_1�h�!Q����� �BM>r�����j�p�|Pr�rZ=�M��9�;Jq���2�5����*c�7�`�@H}8k5;��@_
e��h�SY6/B~B��QN&
b���I�[���Z����3")(�[*0]\P� ��=Sf!
�i�qg)	�Z���v��X�$�O�P h?8� Y�əe)~�Z� {��"�w��0�+H����2)@��Ow��R�\Q�Ղ�_G�	���gi�Б	��J&�"�-$[���k���Q�(��`�
��x��Y��P��ЂIڳ�b��|����>Sk�$Y�Q�@%�����]1']"�Cc[}$ �FA:���*&� t]IJh�'��4�|��s���EY�l@�K�D���X�.������/m�QD���-d��݆�z�l�Dh(�r���(��]���`T��v<?�jAcCe�zzG�x�4'ћ�h�����7.��<B�� ��
�z ,��<��OF@56��]��z�L�h	�2y��X�R9�u��`;�9aja�p�w�][��YO�)݇;��-v���Y+vj��Zu �Q�K
p�ډ���ahnw:����� F���WH�%�����p��'W���b�k%�|�,R�@��Q]e��kga��/A9T�O ��&b	:�AI�h�%pZ]Wc���r}^���Ԯ (�^�-��.��-�Z
��#;V9'��`i�9�&�v��@�Ʃ�P���XV�����=d�3��w��-T�K��s��Tvb��CFt��'A�]�'J����<L�dŋ��oAJ:��*�i@�euph!�[ ���1��MI��A���<�&[���45�X��>��p/�f<�'uÀ�! Z*e���F�	]��O	ށi4 Uh#
�Zo��k���k�z\S� �L�D%�t�o�_J&Up���L�AW�k	q� 5�lY��Y�rމ->��LT_�9)ʪi��O(D:�������K�Y-<��.���"6s\RU��>*��~%P�cԻ�H1*8G��i�'_���;�J`�K����ǩz�AG}�А�O"�3;Wܮ�q ���URh�6`!*O�sWD��r [�݂�(1Ŏ�"h�e�RJ��'|'[&n	.��l)%�����k�����8>g^$[���p�~X-k�8ţ�)G6ȋ�N� YH%;i�{4/gM!��&A֥>[�B�^�B���6�� DB,(�-�# fRQ��S�������{�������p��h%�X��L���������j�RjX��t��Dؚ	�_ e��CM$�2I�"�7A��Yu6������oKՔFD|��ǫ���1s�'�d��XQƄ`�ILֱ�U�(��A�! f�N.���/)�(A�BX4�!�e~�c""]]���1r�-A�*�^>�~6�����Y1Jk���ZcȚ�6xD��{����hKP�Z�1�^aE],/����@��e��}�)�Q(k}hf+>b07`(n^�ʿC��PK�X\'	�Z%�����%�8_�� �@D|;
]��'�u���|����.���IR|z> G�w��C���I�d`�í�N�w���#��/@ f��Z-�`�cv ��g�m�����4W�P���@��]h��� (9��J�s$����Wh��tVb5�	�7�(���Dn$M���� �v�x�y_0Yr��ֺKs�м� (�����>�ÒʷA�"E:)�T*a�g�S�� �NDnl�x�-��������Y�v��Bm}ۓ������/=�?J1B�^���n�"�����]���� �j��yT�A�.�~�f!��	T��=�+��;���~sQ�,P�aU:��n���X#Iպ@����2��D���!M	��U�u�KUS��h�U��z�Ш�_�HOa���5xn���`e2~�KP�� �>�����z	�T$��P��Xq �N�����qhZ�����4�@��Y\���+���X��B��R�T��`�S���)� ��%,. �:<3�=��	�[�q�$�?NK�I*I�	���m"�Օw��3I��P^�GG	�Ax�,�nt�{�%_Q�I���q���v��>m�F.-c`�\�G\�J�@��@��Ǿ{�ݱ����S+?l�!3�V$ 1�^C�keF�
� ��h��J�_�o@�)J�KS�c�*�=�
�0�P�1^�4�?@�$@,.c�(�� 1� �F ��1>� �ی��\bE��7�1Qk�gc�(�J��0�d�y��1�se�Aё�Q1� �mB.@���qM؂c��~�I�!��������[N� T��wfiS� � P�7V��)\1�Y�+ �G �Mu��@7؈N��)H؀�����������;�g�@S��@��@��� �e���� ���7r
���]�(a�����9�s��&��,YU�P��Sܣ����w��j���̑�t�I��D���Q��GR����R�K��/�#��ҹ
@����@{bB����@�h�>~U�5y�s�o���h �� ��c�1�*cq	��10qic����@��d1i/�9�@#�Xb��<�ۘ$(�u��r�9�D|iGk�( ��I�p��2l�Գ����8yH|�=��2��h�CX0�m`���ɤ:񖲆&��O��;G,u�����=� D�@I�u�,�t�:� Ѩ3���2O0,�]�XQ���^2B1ߠʳ_�/�^c[��84h%>������9���NR�-9pS`��
E3���ŰH�2�Vǣ�w8�>���Z�`�8ĮX��B;�u����PJ�`�+ �	8�Vp�bKJ�傞[��(�1'CpU%��~q����Z�?��}K��3�)�3�XXH(Ϥg\	Y��h+��A�x�u2�tj�M��j����N��of��(i\K�}u��-H�jr5�p$:PH�l��$�EY�X)��jdY��fK�����ʤ	��5Պ�Y��rdu�jI�b�f�D�@��(�Gp�K+|E��	h��0�gG/�z 5d�.�7�{ S��W�1��0���냦��E �5p|/�}����ω���U��/��-pp/ԐQ�L�� 5}wRWh3M&�^ �2zve�0�E2�,n�O"���1��}D\�b21����_ R�%-���DT������:V��^j�����9F��gi��bd\c�D��s��"�Vk)�Qh*L9�%�_f>���2m2����(}�4`��V-�	����0��-ڛƟ�z�!�]{�n�h�|�Q�*�^�݇�P�Գ�X�Za'Uh���#��h :j%U^°f	�D���K�@���E)��7]�0-����?/�3ti	����|�+1�6�Ը��
k�[@�4rp S�P�y������y�:P��(����uP����%L���|��X[+�y|@0�鲵�����=H:}� �W�vG�f>���3F|�^�n������J���R.����I̹)G�k���v`pA�۱z�Ap�l�O(�O�,
��J8ưk*TC��f@y� Y�g��LO3�wN>Op�^�������K�M3�@�2� ��x-L��� �����
�h`��3�{LccQ��s��K"	�9�p0j6 ΃
���\����.)Y-h�Q�k���p�~@��w�%r]v��suM-����h�^���|�}ﻩ&��&3�i%���JHF
[�4)���f��8H�hI� ?�/Ov��4�q��0 u.x���\f�!uY�b���������t�h_�n���T
+�V��3�h�7�%T]o�*�����Al Rh|=�b��#�q�lu$�p��6ǻ.�D~Q�)N����Ȣ�(P�]`qo�2�5K_���I1�f$�A�n�:t�1[	U~�h�A�`Ng^��J05(�B�h����j�:	���b�3�r�c?"z -5%I靘e�Y!��Δ~�vx��Q�MpnIJ��Q���~�`#�m�n𮨀�.T�hE�pgIz�\<�U �_zb$R
A�V�����̺RYAqU�؈kco)T�,����h�8Q.�^�&e��.�S��ShH\�n��7�J�g��o�w�k%�/�eM_qRGs_ӺEX���7>�Z�	h�/;J�MTj-j;��(�@�﮸�
)��h�Pم��Ы\��!S-z]h�~��j��0�h�B�[䉊-BE�T��v@G����v<B�y�p�MY���F��'Z(Z,�~��r�2U�8_��|u�+��:���ӟp�|Ԛ]߁ϡ��OA@��.�K��d�oOƞ�ZXv�h�#1�A��� �gǛ+S�oj҉h�pbs�&�	5QR	�f�ń鮤x� ��Vh=/�^����$��@��Tt/\Z~�r(�+>0ƀ�⠕fX9,�?%�D��X!��#����x�]H�=hλ!xR�n�����i:��.W>$C�JA	�Z~]Oc|��aD�p�,k�).�j"d���s�C���%�P�riP)�;�1�<~EN�铤�	�eR�^f-�2��h�T[b���}@l���#�x�����R�n������Xw��p�@�B�(J�,�~�5�"*)�2!�z�R��Hp�����d_�+�$����2�ҙ��@���#EH�����=�x�	y)i�qz�O�a����~�VWN	c�[1�?�����QcI�),����µ0�Zc�C8� �[R4��$�,�B��!��<�"	�xfi��'lW}QH;SG��\��S�+DP	��|!�!(���8��[�} -q�bX�"ʾU	>'&]hn ����xs	IM� V��x��OLw��D�!}�x.���]�\�$���/�����sL����MQ��n�Ϋ�)��_0|%F�Gq�X����|k�5\����n�w�&w�����)�գ̌�_������l�$I�j ��' ��c����B�m��x�����@NEJ��s(�X�:�qh8�uTxH�ٸ,
hE2�i��o'�������814���л�k!����sT]�Bx7���df�F�I��n�28<dpT����or�+.N&�%sdV��fa��Q�P�優��4��,�a��M�n���b	�#�j�T?��P?�^�yh$�)q|r��Phoi���9[P��|Q`l'L�r���h�"�,^ڷS �M h���\�7����5'q:ak��-,���g������Q��S�H0��������(K�a ��Yk��/Z�y?�y�9�P'
��H�k	����q����&-+�2R��HX������^-��8w�~p;�Y�{��h�L��c��q"=�/]x%%��]4i� �2F�-S ��j�%� ,�A�5="^��Tr��4T��-�%.���9�P��ݙ��ܷo�I����� 8�u��3���'���/�M
�!O�Vw�|�n'��r5�l`�#&�GҬ�&�� �r-2�[Ѵ�w,n՛d^�C���Ӓ���f���.��qv(љ�"^����?�GE�8=إXB�1� Up@y�WZ#����@�Z-�%]/7@�+$�K"�MX�ĵg�c	͜�R�"jBI��wF��Y5����_;��X� �iZW�|MlX�\-hE/������_b<Y2�!�Ȭ���nU%�]}�g4�`a�|�WrN\��_�)�����It`�m?@��/��~]���g#��,�����R]���~��/���w��� �2'���a[.$}�!iH?�[^��TPW=F6�n�`����j�X�_ĸ��I��32�,Q(�/����g*��I��_��&�k�������4@'h���
�C�!��!�hLy6�f3�Q�;\�N-��H�N{�����Ӟz��a�
�o��K�%�染=٨����Ú~����qt��7��}�"3�/	��P �C�Sp����Z@�x\	��ۊ�O����q�Ao0��d�G��F;�4��0%n4z�3��@:/_�qL�fX|8���;7<B��S���0c:�{@k: ����-��	�\؁�S!C���Q���[���:��R�!j��B�!J�4��
�mi`���"~���Y�VUB�b��hr:�Z�8`xn�P�A�h�;�y�5�r��"�����.-���u�龺�X�9�.���G�e�W/�N�"! +������M8^�m�(��PB����*�8r�j91�2�PwQ�K�F�2�g�/L�4��
�e��&;��Q*�v��^R�@*�ͪ�(W��T����:d�f�e_�����\hq��0/w��(SD�K�(��N�a�W1�,v�(wJ��jA� 4�~2P@��+Ch�#ta��Q�b�f�;�L*?��6���F���wR�2�����9�t��z(Eg�w�q~�|h�Ss�K��Ks�	�^_�JX:5H�������j�P�1!e$������ߝ�LC'�V�i�'=��W��'�p~��KdO%���\2�9��N�����u@��%G�@�LT$�U Z��}�M��oWF��n&��`Sh	<*|j�V�؅$(���BM�|��� �r�NaZ?h�`3zJ�*T�eS'�0$�=��f.hm�^�q\0oA�J'����	���+Y{�Y��_ ��&�?Ձ6K���;�v�@��2���>��s����RQ��]� |� f�"K����Q�^O������_K� ���0Y%4sK����Wu)�� ���Z|�,?M�E��S�Wa]����zX��ŏ,�p%<��Li�`����hJO�ʴ\р	頾�q��`v�Qb�̈���]V��rk��}O/��$�� ���4�,��H vJ���T��ڀ�:S&O�s�F��rT��h/vWt��O�H��+=d���uQ��5BTb(�)�+�U����
b�=o��>KS{�._�qc��ꛟK��ЖI�J$����ZcKY��V�{��c�(�U�PL��x��b���x�	~N���f^h$W):��[�*����OI�
�C,�A�|Y����7 )M@<�ΡQ� �Y0���$���b���(�ћ�1��DX2�a|*;A�xU�V ��|T5�����=��!�3���	h�a�d��\N�<���)�� mJ�Rո��N(�bVB��s�X:,���3+(��`��0��;������I�lt$��n0!T*�J�RF ͳMj!�( 
7_X�+1Z��,�BNu �/}L �Kڪ\=�H�#��l�O���G��?��������_�[�c�1��.��JY�;`�0]U0�2�I����_HX��3f�$WhV��=����3`��}�%gw��hLOy�Q����Y�[��,A~మI_��`���\^`�QE�6�uW� 	�0��Ɓ�j-$>����+'U)����,�s��W5̇R8h0V� �aI�[���� 5m�U��~��D\���K_d�2�]Fv�I>�"0^�g�#�u�E�]O �Wf��$�� @#�%1��
�^�E��R8����uN��	y� �X�ob*�,���t ��L(�[�^S�	��Ѱ,�%����s@t^K)$��I*�?}D ��vF*��(�_OZ�q�[���^�^���`_� �7L[�h�k)��]�Ps�zJ'�YS���#*'��[��Os��\�����It�[Q�L��.m�:�z�ծ�7	��FP��x]:���M
A��`�xB���']���+�($� �Ht|��*"y�0�N�)!$!1���?�������EPkR���rr�Y�$�2�Z܏P��$�ƑEm�w8�r������B8sO�81�,iש7���*��'ph#�^tXZ��z��C���	��]q�\�`�WAw ���^����^��.S�,�)�Uǅ�\�=�,օ�=���+OT0��Fn���I��R�@҇w�Z�thkS��Q	���}��A�^?4���Y�ϘvpZ�������� f_%T^0��.}lC钇V�=N��+����ލ�2Y߱ټ>��)��o^A�0���[lR	�q��z�(��D��@�Y��!z�RUA�*�G����$��lU����[؀i'�t �{!���	�9+A���#�B{���z�|4I��-'Ⱥ�:,�=��r?�%��1��SwB�A�)�R�P�{�����O��jzF �? =���i0�M0��@^⽀�XN9�(�/�U�.�6$d'֗�h ]S�~�
��0��v��O�V�� ����pn��{����8�[%K̍/�UT\P,���BQ$PR���h*i�_� ��Z'J4��Wi�z��X~^/�@�����Z(�;�D��B3J�ݩ���Y,?܁���`a\{C%����-{\,� vh�2%}� ���Tr�X��6' �������c�	�}�烾�1�Np����Q;�v�� ��('i�	P��xx���.������n�^�e�G�2A&�(� >9�U�KB�����*�Y��Wh�y�s�LXG�0Y�l`Q}�@mR��N)���O+4����_!޸5t1|� 뻏ik�ޝ�,��\� ��/����y��S(���X�����m�H�Dt�SG0� ���~?�Fʀ�2w�M�3��Znf�h�(*d���UQ������	J�'Po!�s{X,u�T�Ʈ?7![����L/������T�%������V�
Z��@#�!���>�]F��� �lb�twg�(�W�&(����ؘ���w�'ܕ�#X%y�a�����'�Z��Y�����_O���wriGB��n����Q�KTk�o�Ε+�@Z���5������'F���=	3eX����Vu�-�>�x_Qt3�k���XL�WW�G�S}Q�D��ü����� �%F@ʼUi|%_�	JRA_Z��7��g����[k����(������tS���$�ٛ��ξ �E���VDU$1f�FP���VL�^-�6g
���&��]�R{���OV���!�-v|�8��>I��K��o�4|:k��� E���{JJ��h�r��]|�,b�ϛ'��� ���-�{|O����C��8i�7�%[�����^���'!�d��)A�A\��C�U�i�� lvz)�-V	�Fw�?��r�%ݷ�wH��gN��q@�5	�:}u�~ւPpm��1.8`����! @,]����V�h)P�W],�W l�8,�	�� �:��1�"�&V�5�@X4VR���z�:�_�f¾V]���)%���/H�s�}hI�!�b�xvu�
h�d��P�x�At�ݖ���3�%F_�^�Ͼg�4�z�kG�F���م`2���c�~���,J���BnyJ�+���cK �Y5>g��\��w�m�{$h&�n���WQ���kz��� V�?=K�T~(h�W E�\�J-Y2��h����{ف�|m�JI�S���ؿd�.d��G�2=���߉Ā�8Ԙ���;����2<��6�/RYѩb�Q�hV_�yK̙����1��"q(!�Ć�����pӹ�� ������Z�yB�| &EN���	�sm��k��X���IH����:���j@ϺI�����^�G��B�I�h St�~�J���v��ն�L�?��U��?��Ѝ4�(��2\��Ys����2$P����]��R�Q�O��,b�m0 Y[W��"F8w�1ݮ�>�kf�4��tRY6@Qh�"�wY�r���G�01�g���&Z��:��&���S;��!��"��Ta�E�"��%fB�6����d=��y-_S�V�I1_���RQ��[�_�[�EGq[�i�? t����sz{��a�P�����EŦ�e03�=���5C�w�������������	�`�	8=�J��˘��Z�5��6��p�/�W�t� ��M�R�J���X?��E0��T��v�,K7\�L�l�E����L4�	kiPDv�[v�o�+�E~i�(5c�͉l9�yA� s�-P���l3��s�C�LJD-�RJ�E���K�'�'t@����un X��yP.1� 9�̈́�	ނZIPӼ�T����Z�s� ����$.�p`��N����i�l�&�'x­kL�}4�{×ھ؞����
o�0�O@�� ��)�h1�w��+/���S��0�(�ZC0�=�\;�\,2����[MH�	P8c=I�S:�~������T��h%[���_��$Ã��:����g�(9~�����K'L�4��~������S\�V��U(|�%�,#y3X�V��+��}P�d��8,vH�)���
�*�� ��M=�p|J��೻�[l8���C��d�$�e���.sZz��?P_�מ�-�dp�@�	�#�Y���g8���J�V���M��3�ŕ��h�^��f6�mN^�f'�_,�H!��J�T���pH��\aU�d�e��S���
I�U1�z�u_)�>�^<1�'�Z��#[+9���@��wfz	�������eРh��IR_0�P� �ܘe*|�Δ�?����N=H��A�P/�����3+�6�nd�1^Ӿ-*�_[���� A�K�<�k �����Q	�:�V�rT���?s:���	�z�d5�v M����	�[ ��W�g��oͽE0G�;�!�@�©�%x5���ÀHYD-�6���=�?����-)�^�"o�]%��v��fе(�m*����~\�-�=�[�,� ��/YE���.�`��U���� &�P��G���A1�!�,� Q���������A`40w�'�3V���a�	����-^��{T�,��B5L�Oť�T��KA=N��NS)����L�y~J�`��'X	�ez�P��G@�60�J� � LZs���������r����-
W�#�!��d9A���'/�v�r�_0k8�Ƨ�S!��S�4����*�_�	�t�-a^�/!�+�����Cc?2
Bh	wZԼzJ3 �Z�r��	�S7,u�g`Jh�VL��X�t���8�vO��	/�C%zw	��T|�.�a�%ޚ�w��$��@�8��^���jT}�_NҨ��\��U����n�%�X��h ��vK'�1H��+F�t>O��5=�q�ʋ�[S4N��<�)�^Z���.�3�HB*�_a��~T9�45Ԁ��!/'A�ÿv�l��`P�&.���R�����/*[ ��.�0j,4��W���+�Z� ~h��F�[��/A�����6u�07�/��A،: �.z�&������~<��8��	k�� �P!$bG~/�2 ���W�^R�O���
H�$u��)��<�[�)� ���E���;�h��ܲ�2[��U��Iȅ�vp��s*Y���hP?�Eg	���ۿ���_�&���*�3�(��~(���QK�� hd�A1ޘ�@X��{����į�I�|H/	D�u B�kݿ)�[��sT���xR%�ܐd����YR!�0�'����b�=E|=�����ү�UQ��{��o4�j�a�y�k?@��	Ttv��4�%�e����yc�&Y`��h���0IJ���L�)>>�sI�mQ�%��}��}6��8[" �_ř=N�͝���� �W0�.N��; �Z�\V
:�-> "m]h��V}L�.��Q�*w;�?�f�b�HѮ�$��u�4ϊ+p�<Y,��
�/�H*ɿ�v��/GB���w���c�fa�6j��+ѿ�~���n���9��QT�-+�� Phj�X �cSrH-�;k�J��8 �e�h7M&��a�{`pnx�p6-c
�N)�� �U��淰'�0O^�H顖`-�1WKT�W4l^E����AL�G�i�`5�S~Tc`���8k`8��̽���s���"�D�^PM$)ǁ	�jB�D=��U�����a�S�Q*�����%C���	hLw4�N,���f��u�	4�0Ƃ��Z~i��ҥeܔ���=��!'���-p<]��4�0�X�ʣp[M��|�ݓF�7Q]G/}�cͽ~�RY�_��?0Э��gq�8,��T:����V)��n��	soB~ en��`�S�O1�>(��i/�*eb��Oð \���R��gBoaQS5�P����.�j((���R�b�0��Ϊ4�^=�r	��v%��iy�Q�9�OV�>�%-��\<$ H�CP�n���N���Ɯ��\rXQQ�~�)?,K�g�N���2+䜝KyS5$�,�df�5�`۽�kH�{EA�..���5�p�h�<Ĳ����:�Bk��J���4dY]����_����(��I5%e��_����n�:��T;Ix�ݥo}�����N[� o��������x۾s�U�;�*R\m���|�{EWh�_)����7w��/n1 ���Q�-���0�Y���'��r"�n��I���v�L���#�b�w���AKQ<H�^�8�dV��#���x;yx�&�w@�9h.E!�.`����Kj�#�'Ši�q������ټ���gu��	*�O���_�\Fk)d��)�P;�^�m��0��Gl')��?V�K�'8 @�u%4m7��8t!��+�e�f�K�`��D��;�c�Ή��=�ZR��y�ч�lNN~S�P��W��Q�+��""^F��(A�Hv@Zm��FD	��{��"��QR��!�*�U\�v�RP�`;�f�"�r@���٨(EC<�}�Jtv��
�	.b���wD`'�,E/H�8��e-� _��Er ��=�C����s �r�Z��ue�u���P[DG�T^U�H8�'�D�
��_^`�R�I(�Z�?e,2�g����6���� %��Q
-X1�"�b�Z�����O�!�����ь;�"��5�k=o�����uC��_��'�Z"���
d+JX���z�[���X�.���A�E��!���/ȝSj�^-
��h'=4���WnzAn'����~���N��˙|M K9h-|�R�B4ZU�W�V����Ů`�KZ�›�a5#�� �g1�Y�IwjHvx��/�Hҫ�e `ԛ�+id���C'	���㒛�m�K� �`��ECc1�I�{�_	���v�Ũ�N�9o?���w��F��0Y��e˭q$��T~U�}I��h,�r��^l-:ҺLW��/.�q�$�ڮ��h�p|7ď�<]֩Y;~	�y|>����!s�k��=:J��ï��2��p�vT'��]�_Q�?.YH�\��w����m�{`w����6ns{�e��K��:kf�1�6}p�K7����Z|ф!6	Y�ly~)��`�[�(����8J`U��������A������@r�5`Vf,W����{	�u�����o�x����@�`U��h-�f! I�'1�}�@�O7#�@�+���_h{)F�݂�Zu@�<�(�wQ�.��a��� YQ�� Ȏ>N?���������(��u۶~r r�
��s5�HLU}I�J��#>��KcE]�����,��H��t�����(�)r�D��Zͤp�E �d�8<Cq�o�{��/s�>���C~��Fv�%��oJ.p]YB�U�X+�t�"3�8Zp�� ����Q��C�-E�N��a X)�Ӹ�o�]>�D�W϶��n��#A�Sx�=1�aĪ��b�y�K�1h*Siw��'`�|H{��3k>��FYb��Z��H4[1Z|�U�����Vt�k��|�K�4��	h�g�,��O�E�am�� 08�BK���gbẆd��y7ǚ����	Ph&��1�����FS�Pp"�\w�FI�mRR�{Pk�>)����w&erΫ040����,t��vh6lVf&���0%ԾݏI�j!P)��ρϺ�(Nr����Y�[,��O��秿��)��P�
�^ᑯ�K�U܄V5�ʄ슔^ ��hz·s�A��o�A���� z����HE�y�G�I=�h߷Nc{G����p�I���'�y�o��@ ��-.ڰ8X1κה'��Ǜ��xL�J�}�=C���Uh��,��cA\7�+���)��/��ꘄ@�9�0 x��RB3���]�o��}����6�:��9f��\�WH�`�-#^�[R���4��I�)K(:�����6"Rf�(N��)\�z_�'���F+h�xJl��[�~q,� Qw@^<)�|'Yf?lP�j��C��W��ZR���`=��5
��ܳ0�,@C��H��b�<P'�3�_�0!�	�)�� ��rA	�=����Q�^#�]�d��+��;=|D�c�I�/�[�>�k�
����nY84���q-����
���@=pij��nk`���	Ѡ~�:�W��Bhr~�^ �)�GXQ-o�z������5>wJ���1�j�L�0���)&�7~=�V�<��t��h�I	T*�����ʐ��(@�A!��{Jj�����D�К�ig&鋡;�:n!�h;�>1ȐTJ����9jH���D��>9~Yh�O�afF1�H7�E�0���m�,�ʟ�[H�ғRA�'"�Pe��Z%1E�_%���J7d�P0��[K|B��q�Ű\Q���d�1�� yՕ`�" '=�d�Eޯ3/��^�	?w��*��H������EƋ��Rկ���W�P��d�[��Z�J��
�^�izH�k�D���)}��x^J� S��w�F����B)���(��	." � H-P�-���ގ1�ɦ�/���f��������=u2"��3�I�-�VR�@_� ^~4?�TEz�e�2�Ǐ�9���]���?�&W:?���	�`T$��jf{|4 Vv���� ����.�>����T˹�a.�uX�+��*'�]�N_PҸ��~{!�An�rV�H.5(&��`�-b�$6�v���
B
�<ߟ [)�
`W���JqJu�e ѱ���%��~�]�`V�T%����ŋ��Q�ּD�P�Bm�bPqE(:� h�	/��l�[�?�5Ҭ�C���/���(�Y��=6*�=�.ي��D��ּH�l*z4 hߖ*������	
g�G5��~�#;�@�Y�9a��d�µ�rx�u�Y���#�����,c�p?��b'���\��
w<���:�_�����(��58�/O6�^qC�Aao���b�.+�d� G Y�0O��g�MC:H=�w��N	��8�9v�3�D��jJ�R����aU_�On_�F&����wKb���E-V� w�	DA;O)LiAB2I���Ηx�v�;!I���\*����b2u�C���OV7	E���L��gKus�،���z�Y��D�or2HT/'��ϛQ'lUG+:�&���%�V�/�Z�Jjoл�����]0��=|�O�{��J��rw�L: r���?��[̑�/�����j{~|z]�@?�	����u��(��=NBg������^Y}�N�9rJ�O/�5��Q��S~c�T �RW�Vx�&x������wZ�Y��HK���}�D��`�d�d�"�� ��4���q���(X�$u��0�7ݰ5+)"��z��:1r}�A��~b��)�ཇ1�@օ�+���&K-	�1t�X3_�H^�h�K�}�
�5$"S��`��+�ҷ<'����'�͌�'z��H�$І�!��Ӛ�ф�è������.#��^PZRVS�Xn�(|9D�h����%�Q)�-�<�(N�ItJ�+�JX����V}!���c|�1�[;�TԎ���I�e̄�&"|3� �����-O�,�gk~-�utF�H��
��pk�1�L�����)��IOi$D�p���9�U�D��/MW��a�� �Znj�+%]_塭��r`����e$}/F��v�L�w�[X�.�e-�]z
N�(�8����<��A����)�Ѳ��_/�I�U �>��7�^��G+Wf��o��Y[��5iE2�� `y�)@�_^Q�i���S0ְ_��n~���\����'�m�Nb����9X�=��`C����UYQ$	����M?�R�^�X�yNx@NY%:�����Kw���S��]���'P���<baa��2� 
[@�w�Z�E޾D3�W�2����9��%A쑒�X��)5OS@�Fj��N1�X�#�\] ��B�Q�]-�_h3o�`��m陊�П��,�c` �i�^����n�P��Z!=A���Oρ�<��x�F��YN�Oj㉭	}�g�f-j9��tW��X���Տ���1�L^��Z=h>���@DV�N`�sFS �] $8�$E��uk��T]�.�ONK��)O��o�0��	d@���"~��},,pյ��n���/����h�@[_*�� �i~���k��Vd|hJf�����w�!�_NjB53wpp|'�H��	�.��C�
��0�@l��`��c �S��~�����-�_��$�@-Уn�iJ��C}4q��Z�A?&_�-��n�X�o�Nk]�[%�}l���g�`�[�
�èJ"�ˍ9�%hRW�A%	D�4t�_A"�2�Ә����[xH U�!'	hN��u^����	�+��JƛYŀ�JX����w�E�b��˳W�[i u�}�U-� ye�J@%�<��0���uS�@�`bak�?�h�pcH��i����	Eީ�Q� �Yvk|�UV��5�^��o�X����A�,�rC,�uX�i�:�^�t���K'��l�k�՚O�;�>����k�  ������pSwѐ�I�.
	�ǮA�a\h�N7�U%�R4]��x����37��� �-UxK%e$M�q{]5��O ��wS'1�|wɀ��!B��['TbG��ubKzi��Z��T^��漕A�[:����5�����2n�,c8�ߖ��7K��΄���!��,$�SH*T�ܣ���R��n-p�k1���	�+ �2��Z!�����<v���-������襱��80;'A�:�/�ay#�Iγ�x��	�O�3�A0EKD�� S�c9dXK���E���"�@��|B��M�����&��(�J��q�]z������i�0%�V������/n�-��.�<0P�#Rw��G��[N��ԫp�hyr�)�1\	+_Gq�f�L����<N���t�@�_7J�:ׯ�
P%�����隂&5_@��-xd\5�T�&�LR>A�'�^�=�&!QS��-v(4v|W�D24�h�bF��(PK���(D���`Z\LJ��	X@�1V7��IBd�c�-�f�i�>�]R肀�0U��� ]Є�h6y���Y�9\-bx�K���	7gR�� �$�IY!W��J�	�Z~F,z�-f.�ɭ&옼�Db6R�8�r�,��H-�F��	h !���{�������wR������_����`89.R��.�6��&��t
�G�7Y��]喰��YEJ)��'��d_B�_q�k"h��W24Z�.o};�4���Rlg����JT��OM�h@��=g�X�����J��	U�x<L_	}]\Ӎm�.�t���a����	�F7����t���1&�-%A�����	�}�B�i�?�Ѐ ?�ח�r�/����pe���"�L�fd�g��7*_�܀y��<e� ��I\�#�D�/��Z��8��jt���[*�B0�w����p5�X���K�'|��J�K�i�]Đ������ߜ����[^�d,����  W�ܤS�}���Z����IUmsM;c]uz�<x%�w��i�q]z.OY�2�Z�LhN=P:���R�h=B��C��c�3�B�s�ة���.�P�lRh�3-q�LQJa&�Gn+y,�Ʈ䖔��K�#!^P�<�]\-�jۄ^�VI�����`�c/�|a ��M�^W X��gonkU2�vE�t�B�3Y����$ʞ:�i�ݱ�[*�URB�":;3��-�TQReR�O+�u��}g�m"�'AD�U����%l����{/��!P�qyan����N�HPV�ʀ��#�T	�����̷�E.&��4��O�X�0��?�[Ӆg��S�{�4Q�,��?^��U��+���A(jq.!�(B�����l���\�9�j�CX..�11����;�fH&�n���D	'84R�8��_�8�h$@U$��� -�yA�!����=�q_��C�E�s�r��:ʲA%_!���*Ʊ���EyS%	��Q�Hw�fs�y�*UE��Ŗ��k���2�HSX�=��W�?��	-?�x��<�8\��	 ����в�15������@}��U��[��ofŰH]���2
B��o��h�-V_��Rī���S>���s]&�0b˲��H��	1��I^i����ZU�BbP�STޫ`:�O%)�gሪ�<��|�B���oI&^�I�}�շ��v��.��*�^j8Հr��LWlT��K�Yu3��D�v��y1�RS`�z��%ZJ�D�
j ā�v^//��h�1
`8|O 5�k�b���� X[D>�fh�Z*�����94A���昪eWԴ�۞��	���*#x�������LꝀ&2b9���0�����o�_F5������� |Ro%����[;������'{����Vʤ����P^��1>��X��������Z|^K�*�J{QM��,%����	/��%�yX��[(���JY,o�SBhG@�/���:��{�S#��x��^��X���Pu�i� �e1�<�^~�a2�M�0�M����.�S=>��*�C�Nf;H�1���k��2W$�Z<^���-�.��H�x��@`B[��GUg,��8��w�,�4vA�zr?V�av+����\K2k-���:%]���ޭXw��;��f���6�*{��+�e�������N��Jݒ�(�0��b޲���9:�'��/,l�6��[�2�ܽ�a$5H�]�Z���J�,��0zqf�Zt	1�] -�d��A�c�J}�a�G|x�
#B[�U|>��j�ŽRV�X��+� S��@M���'YA�3 �h_rV��~��� ��B�ԑ���퟼���TKX��فώo;s��;q��{��[�P�[��O0Y��Ѷ���d�-�s'Lx�	���	�Rh�:�%���`+��BA���i��}ZǓ����hS)�[�s�;�4K�亅΂�(_'W�ȥW><V�~0�P� �	�n��5I�%���PV�����]40 ����0��B/�H�8L�/�f�}H���h��5�,�Z�5a�B.1@N3��;%We7����df�~Z/���h^p3�Wؐɞ�m��`#��Ύ�	��#�@�HG�-���SG��d�%wo�&����%�[�Q &yvPJf�"�$I���UX����V%�<(Y���[�XxǗ�/������n	�����.�["�$e\��ڣ��_Ao?��� �;1�� ��ˏ�2�)�Q~kX��x��b����"K�l2��7=�/�XpX9���X�	PWE��_�ט�	��$�id��<@�Q�8���]�Q��=|?��Y���� �9'�ĽTK�c �H&(�p��Z�Ę�B����hv���5V���4_���jS���w�n��Ҿ�
�.��H,R��L�c� N5������*�S	��{o\��}�HwjJ���`ʫ5��.�R����Zp�:�,QS���΀�:�ѝ��UcJ*�q�{�Ip���y '�A�n'�L�bWgA�]H|b0v�/9�rc{V���]�U���~.n���rh�5���W^E/�7R�V�;_��� Qh�H�YޱI;[vzp&YYP����ϵ�������_n��_���yScр6W�`��-P��)���U7�p;!	�ȝ�[�e0W�7�na�s�ׄ�(��������=%�<	���� �YShz���%�g��@e:j,:(���%.4k��~�Z�	� ��NL�]/��P���g0��R��{��<,s��D �/�^-	[jC ��A�>2Ȥ�z	1	W������N}����[��j�J���j0<�Y��(�,>����wx~0@Ą�L�@��JB��J���e�b �^�o��s�,�"u-��P�Q��uFMT��)�ԀbDZ��1�Y9�_DƂ�lുKWSV����ٷN!�N��8M؎ŕVSH*;ఆ�q�X]�S����{�����r'ǩ�+��r]��	��lA�����B�<�ـW�R`���%�0\����"fI y꘨��1&0'hSP?�7�t��z��0�v�Z� �ot���-�R� �@$X#�[a�މ �y'	��_Z��i�1���k�&�Y�p�ה_��%����VUhZ�E`I��xYY�뤭�)}͕�/}Da�2oa���_�]�"^�B _Rf��>�n�XK���F�^X�ꀜ����](� ��H���5�j-Ĕo	�!�@ey#-�s�Bb����]�l��q�54.�K)���ZH�_�J [� Y��6J�	I����~���Q)��准S�������� �4��RPh�X4�%W~85�Ĵ�;���Eۡ�{uI����D7G���\�Āʜ�Xw��~*�#�@U��h*TR�tO��_�HFЙ%��5	 �z/�Y� �d�����X���*~x�)�VkR���F���׻,?�L�E�0B�u�DKmYg�_�
�Ԙ������VJ;����N��Ug$W\d�P_-�"���uL5{��!/5�`r�[{�@P��I}�P�w� Vo[-g�FK]�Q�Pm�F�#i�-h?t�%�ATwqym{���U�l��a=
VS^��Uo /@��d �s��Sg��/�%Q*,%�;1|�ˋ����	Ý��d��~��[���Z)(��n�W�ӡ��8?�^֊���[(��p�O{�d����r�d]E��l\��s>�{���=���J�F�?�!=�e�N$u��\D�)�r��?2W�%� D�?h7Z���)���ڻd����|��)����[��<������r�3=J:�����P|2�	�B�5����+ʞ��S׭��M�07@��n	)�{AR��fX2`�����!���;�(���ve3��iԂ�¹k�����3��iܱP��Tt�`�鲔�:%}�B�c^�����V��Q3,U٩@4Ile�&��kRh�+A�Ո{B�KUpw �WQ˃�jzԹ�� '	��Y�"Ǖ�����&\%��p�X�*���`� �1�]Q�o(?��	y��/3W"�����8�*+����.S@��>O)�.�/��z��!�t$ "89GC	5�b�(��ࢪ��&%VuZ��O%��� x����"�R*DQ�'Wy_�̨pN�x��L�t����c�F.�3��<�A�����;Sh��,�ɀ�"��ߔN'�W9O00�(@�h	�+Y ��S��
�E����	z�uY�	k�f�(]�" �o��e	�A�`mB��}qE��b,ϬLEf�e@�AP.;$�/��w+"��� ����OO�a�CB[`�#QH*��D]J�� ]��-�K��p��tOru����f.ev� �sX�	h[��K��æD��qqH���5o�0^q1����Eח1d�)p�5	`�%ޥ	 /�ӎ�:��`!(����
��{�Ś.:.�X��[����C�^�� ��IGvK]��E�����T�b�^�}P{���&e�~�N1���������\�s>�:��ܿ j��kW}	��T���{R�`�O�-!@j?7��W�?������`�~�hV_#�aX5,uPH�O�N�m�,�_)�-��F�i�L����^�`�qY
x)a0(�%h�A0ɜ��O��}1MO5�?�� 40Jr��\X� ���F3s�W김�vUO�oPJ��]��UX��LV}L�!Eg�m;k����x�ON�Jb�p �-MdIe�*)�>�+r0��	V����̔.	U������3uY�P�	錇Hh��N_�K�S�D���ݾF�4l9�ZѹJl��ݢ V�YA��ΌN���:e@z�U_���95�V�D}*k��> 7�5�8�F�����_���� �=�U�����	4]u�ɵ��`jf�@c]8;�R�-�K�i�jf�}G�&eXh������ذ7%����C����~E��;���1�٢Z;�j�b�5L�UJ�ϩ��	�u�	Jhj_YV����`]p�/m�*��U�f��|���;���h6�����D��i���#5���H[?��/`�Q��P��R��B��Zr�>�J��ˎO�x����߼(R�Z��H� ^E����>�IJ��횂Z�5��l�h/:��IdaKU�t`�&ŭDˍ�X:�[VW#��б���'WXU�]Q���#]�K�0�t�[ˆ�����&HY���DN!v� ��\\�pl6��Č�Q3{�������f�~�1�[!n�E�
��V�	�^�XZ���h�bn�w X5�O!׽![�*����?�R���YC�X��)~ ��] ��BZ��)�|RA��VT%�����oF}SA�gF�r�b&�N� �6�rK��=��G�������=�cr��S��� c��4A��\�_C*Y=�J�ީ����-�����t�P&y0Y��f��"x	
�%|�`��)#����Y�-�I������\_s	附���/8
%4p��Y$EQ ���i]|Z�{�\��;�zE��Y�+��+FZ�HxJ�����\ M��~J���{��
M��u��L�U��|���i�(��ʬ�]���<k�j�%m� W�����`0�0�Q>kPh�7] �'����&�= &�d:𥲠�9mA1���h�U_c�&Of�8
�����ӓV����QJ���z��%�R���l�,T+H���صU0�2c�n�@c��r�q$���K��4��x���H]��{�%�@���;�q��7���;�g�!!yn�pŲ̺���h����&������qs�Y��.l��cL���@U=�����������?��^�����m���
�a}�x|$s�D�c_�@W�� p�ND,�e����(�|	S�R0�'<�VD�k����0e��Ր@?
c�C�G�?�f�� *�\��t��$hk.�`�����I��^��d�! ��q�a3��w�s�hE=�!e)�.���B�� �s������G)���K�S=�8:ܺ�f[~p���!`8dO�����^�1_jJ{%5["F -,Q~f�I+]]0�e�� �� )=�A�J(r�sj��k^Bp�uP)J�ȝH�f�~A�j�%\}�Jԥ*�;�>}%���e[(�lҲ���K
�������;hT�d<`�φ/�S�'�cx7L�?�P@�hUe���f�/��'�So�k h�W_��*��jB����m��F���D�v��.�����b"}�r?,q���7@�[Z]�#�zpW����=�.	G1�L"�X�ƛc_��#�o<N1e>���Á�,��w6c`X92��!X%��5!�T
�V�d�t3�W<�@�P�:��y����� �v_-\E�&��<)�	����r�0�|]�h����þ���o*���}��]��v��Xs �4��ǥ0]P�H� 8-�*LC���E.�S����y��x`;�t,�Z�a�GX�^ʧ{蒙f�L(�@
[90�0��ֆ���Z�I��$��+�R�R��{;�E��xBO�n��m�������j3�Y/�I>�1r`M���J4=aŽ/n�s�xJ����	1�W>ԣ��{�_g�_�)r0N����/~�#|��,C^8��`4/TA��$:�~	�.)��P��|�5��U�\R�O��yq �6���j�P)Ђz-n�7`��D �.	jU�R��p���k �-c�*鵻���Ho* ���3��'4�Ԥ±�s��WA����0�՞� ��P1Fx��D�T]�<�8l;N[鷄�zS�%F/�_��o�O���w�&Bp|��e�Ҳ���_��s@Ԁ9ɣ��Z��S� ��)�:�ޱD�6�*�"�8x �L֫�)�.�п`�H\N�*$W����\�9���QL��Te�1�SK��L�p�_��+��h-x0N�%c��Z�o_P�$�-�&b=����ok`:U�Q��B�Z* \O[���vX �!z�^��!{�V�������fhd*�Q �ɰ�,(�����^0�q��E'���`�z���đL��>�gkk	'ܵ�-�8�(}��^�%
�"Bk[(V'�,@��j�CK ���E�ڝU��$s.V/	�Y_��NDr��ֻ:N���m�yн�a����~����{���y��S8�
hie@��T���4b�ӯ�' r���O�hc��j8]���J���H��'`�lC*��)�ii��U˺�{�o��o1�_�*�.��͏G/Iv�%�B&���r�K1�?c���=��S 4[M�w�rP�R����0�4��޹ 0S@$��}DV��sE�T]�f�j�1A:I�[�}h�#���Ґ�Ņ���0�w�	sJw@��e�п�Ds@]��I�A�7[_e�%q�	��w�f�!���nُ� (�-<���u��8��_�ӯb��M�P%Zd�+�5���)/�;��Г�� U-%��:4������wA��]��eOZ�2�א��M�l��e悛�{�/��Ṳ�ݚu��z�,�Z�4���*P��Lxǰʢ̜���]Whx_�!��b��k^Q��~�C������?EP{4U_�q��q�'�� c5�=�0�.j��wGl4�Zf�%[E^耿'��1�T�%iZ~�s)���t/� ��GW��D8�X�_�`��n7r��E��p�j�K��H���e����>̿^h���L�M�6� ���7)�J�]�P�̴�ݺM�Y�b�����*'�����!�PU��klq������_�Nt���vq�oyUH�g?�O�H�3e�؎,-�Cf����TY�t�x�Ԩ�t%�1X$sјh��i�Vah�8L�W��@��|.Js����6h�fQ�I_E[���M^�Fi�]yB�(��}��5�:�k���^�!��R�^w��C3pKZ�֪ش�A�/	&]����T%�x3��	k;Dd�θs��&?�b�\^1�S�Yw��fl�����2�YW��X��� �ֿ�`����^�a�T�.蒁�N�0lc4�\�cXY�8h��z�U���h�v7k�ɧ�ؐʲ�Y�K�3��}�l_h*UXB0vǜP%�=_>�m��>G�]U��
�zr�fs@��*8/X�`��D8��;�h��J����KW��a��`:�,���7�q=܌"_®0a�%=��I=�5^�phj�0���5}��'B�� ��&0��eDP��"\O/�8O�1B�&����w]�O.�+!�[��h�KY�c������82��>��NZ�a�BW�,����>$�+%�\�i]��KI�D��Bz��E���0�����)K�%�s�B�<�b�0�4C�ղ�D�C�ߦj��섈⢴��i�\.�M� * �'kʷhr%�$����p�8��8�h,�&�H��M`�8�d㙗b��wZR�rLK<�+��R.�}�4�bFku���e��gA�� _Uh'��*��\�u���!4@�*c?��0�1a�X��^� ��o9^����	|�J�`w�WE�Ẁ%G�����IS��,쫰�󑈗S�wleВ�KG�'�ү�U��yh����[G��r�H~M�h�RHf�߉{'ղ�\E*�hB������aPߔ��j�� �g)%݀�*h0N4� �� �J�f�>)��,^¨��q[�Ð�EXZ���CS<�K~?]��*%t�['LQf�/2e�5�����yl�طXK��zI��%|q٧���*�ޭ2��k�E�0e] ���h�����Z-��U�,j�%u�qX��
��#O (��0��S}��i@�h8H^�r���2�
Z�|]6 4��>UʆK���r�zQXx[���4�� ���V���c�Kg��Qj�WHZzE�R��?O���+j@�i ��!�Y��Q�d���9K��lx?���_d��3'TW��G7-ч�s!j`��J{�^����Ĕ��K�K�$h��^��%a e��7�d�y�$���
l`��mB|&��9�Z���E��»K�K�>�(�UG?�%3r�jכ,��J��jZ�����V�l�����@�"�YX_���! T�3S��[JduA�H֐bDL���^-D�e`�opg��q|��/U�t��UhLl����N����oX�%%X� O��U������"_��Y�Q��{��}��Y�08JO��cuGyn��
h�-;�j��Z��`�.�l�@<X(�T��b���Z�؎��2��lWh*9�y�e���H�h�RF�n�	 �Ժ���,.(���Q�ǀ��V��@��w:OѨ�D{�hl�F��l�I���
,ҩt{.ooe뽭D`��J�~
'��ݲ��p+3gkmHC0�;�d�.!�_�-į��%n�!_+�b��U~
KB�E��"�y�+J�pQ��@�t�@���M�D@�%�_�0!������0����Ÿ��Ox�Nկ-�.�Q�W�Ԫ�7
�N�+t	�> Y��[CZ���	��(�T������N�G��%� ��CD/S��&���0�y�z��6%1뱆`�q)�
� � �?�:��`�b���R�wQw��Ch-yuQ{� �&p�[l�}Ud�()X��^������`y���[�}ߊ�Di a��N6Ꜣ�%U�5 {K]�+2K��[�H��сPWAy.����Gj��N ^7r�
)�-0�h��[�,� "� A�O�fh�G��Wk�T�	�Nk�2:N ��cAn!5.�u���p��	w���*�!�[	��.%c ���1��${7�w�?��̇h��ۏ%|"=��R{h_9�pS����=(�^��O�a�)�*)B�h�t*�����5q-�W1�A��� ���fO�?�A�Y�	:�dVJR�d �x�IhK<�Jb&��`�uY��W�T��~
��cTY��%�q>���6����.7U��]���hps�VTLX���)\���o[�3�d��9v�z/8$���3�/�\d�"|�r��z/������E� �4Qd
�hk�*Hؾ��d���]���./@0w	�W���OKU�������v�^��R����僋��#��ݼ�*�<U�� �%�����  dR�� �����W�<�{��܎0/�FK�^��ҩ��Yh6kz19�>�0�fX`�t��]�/%����\W3F���r� �V/�.~�����9���H��ԣ���?,>Ӆ*[3GVN-�aD���	�A֨/q�K�
�%�l��R2^|���&I��<�Y��u�g�
�6����fk���Uw�ҥRI����p���6��6H��\(O�t�������D��l|/������i���x�:��v@��j�6b�*���Y0�.�7����N&B����>���J���\vĪ�	��JTD��O$ހ��':`U�w����N_�<��[�4��:p��)՟p���W�����[�|ي��@5�3N�S)[��1�����wLk��Z��^;�_�AרX�]���
�l��dea	¥���ΐ�s>�t���/VdU����{7��K�W�9 �Uy����Z��`鹩݅�N5j.�M}EZ���t�%���-ЯU��j�@\����VuJP��v�;�.fP��T��x�'koĹ	_h�-y�	*7���W{R�a��;�ǁ��TC�XB�{���x����S��s����hD�.1)��|c���1ȟ��t�h,/	UY���	��dn�q4�2��%��A(����%,b���5�� ��k\Y�^��z��cP�� uH����� �i=-��.0E>B�P���~����cn0��b��/6���q�R�:B�\m�p��!t$�ei�m\wq� .hK���J(��K�c�Vmh�d��-:Yޒ��mC�.Ob��V�RC�,�̸o��7��$f�	! ��1�`���-X�J3����:��{%K�uk�AHj�5@�
D'9PX�߶�&�"�h���M���ɂ܃_�T �#AGbx��X��� �Q$	�����C@f:,'`@�B��Q���N��f'��4w䃠=C߰)	������[����o�V���py�-2��#�	xyt$zr�h�=%�e�A���+�01@�Xh'�;�������@D=I^Es�SRS�0'Q\GL�Y]Tph�_&1R(Q�u��IW�5#r���a&���]+�W���qa�6�bu��uf�	�=Dt�5��U�B�w>E)�幓�.d�y�.�9m:�wЛe��8�5�����u���,�X{��0�h�Sl�����jY��%�,[ZQ���]A� ���J����x.�Hh�z��O/���s���O��$-P?���#�c+�e9��1�`�IJ� -�A)���	���W�@�u��p��P�������K*/�Hz��bO�Ԙrh���p���K�t���ȓ�0�h�Q����-e ���*�g��_3;��"{y_ aNh����C���G�dc
����2abO��W�pC���[�h"fOiv�x�\���Z���Rv,z�5����gr3��;:!�0Y������Eȃ��l`�ڇH!��s=���p�/��������"6�O;�mZߥ*VB��Z�T<''Ғw��]N�H��\�0I^, ��I:*cM�YD�T�Є�)����'CrST[���cJ��/��� [$���{�je�85���Ѭ��hz['1��|>��[�0�QM���.@H%7;4��3)�QT:��� -.2�xk�z��{��hϋ��%�_�$�wqAa�pPu�ܝ����Twpq�y_Q��>�a��U˸�}f�K��J&h�RN菩 MәĤ��͒�T�lk�Ma���!|j%Xp ����U!�hs 0#�\	��"���X���}�z;�=x�	-�sy�htT^���؏�[��"fR�%vW��`��u���Lr1j ��K�)h� P��`[~:5��)�V���k�z�y��/�+�[Io�\�-����N�/�I��4(���;J}�}�ٺ"-�i�؜K�r�ω4w�Ζ Xph���ҁBؼ��v�G��;�4տ�8�a�/���l��W{�8��ײ}V�I^d%n1�#\
�qh��_43w~� R]���K�kK�"6"��]9������VBE�=^�Z��W4���	EGa���Nh$N,�	�`Q6R�[��;d��Z����[@�$�8�}|g�镐[)��|���K���g �
'KT�([�k�u� �Ә��ߤZ�VAR�� *�vY�?��w�t���]�K hG1�j��Ip�����o��,	X�TN/���%��d{��K��K%[\Z�h)':`m
��z1%�N�ŵ��	�&V�\.�DQ�j�5�:^�=t�^ڒr����w&@i)��@���S�S��n��+�.D	�$m<_��n�(� 
���)�c�_���{9�`��$i%4�U\�Ԇ��;�z�����H��1��ϥ���T�D�tq�R����U�ՕxD����iW��4h�x@��K��<!\�\�xJ���dP�NJ��fW�;.�C���N�,UԅRI�T���M�^w𴹫�+/[��J]�t������g���r�wU�-�o<��'�t)�B�
5 ���(h��@#�X��.h/���Y��y���~�腨��f )y���	S��W˭{U���)��k�JN�D�iW���hZ�Lm��P�6��{��C��ƻ�z��Y@R�+X��B�8[���s��B�3�q[\u*t��-q>�h&�̖��ܒ'���F	h%ȹ�I��v��2�}�GV����R�������h���E8;��>�f\Q�;P)îJ��������=����gkQ���&n]6�MRgc��Aւ���Q%�F-0ٵ
)�X�Ş�����ԉ�D9��΄Z�l�h%8Qf| Zt=���MX����@b*��n����h�
���х	��P�e��h�O����h6���~]gM2K(�� *g��GS���':���ـ����*���5��itWn�;>R"��A~��	���q_�Q<����wfh�H3�L��f1����j�AD�~5��>SGB& @-�j��s�Uʱ]�D+�n{�?+�D�dA\�r�l�@B��9Q��xB[h_CTh��8���O�����f����v��0IP&=(\9Kqb<A���/�v�S1���:�kt��e��N��:�(�ð�k]1$t���' ��3����n��Q�'!5���Ah^f� ��c<���z���L�Ie
(�^��,L�N��ncU!Չ%_��@���_m;�'~�/Sc qz�!�Y��װ���.
f<w�^!�6N�j�c>�@�l�p`X$��d����F����
%F�υ�\�O�RҾ-~`�1(qC� .~��l-�p�Jش��E�m�$��w�o'�"�����ϖ����ff�,�y��#2g?x��꾢������� #t�h�+���e^]�zA(q��G"�BhY,�a�%���l��/� �8HK�z;�#�u���t��l \~�̱j�GRw��r��uVoX8��{��o�|�	`]d
�x�~%7~A�[NIW!�n��Е&$��[���%v&DA_2�4Е�H��t/��,���t����hT�^p6�_6X��I4��>�D�,�!�F i����6���a�q�Y��B'(�x�v��i�`�!K���� ��[D��x&��]X������HU��J�c�XK�Ȼ踨Z��)��g5ד�~�N����p	/XA qLf�۟�r�\~Z-�d5J����P8�T��w0����6=eA'�˵���o[�P	9�ә���^��'/��3�+40���St�aA�i7X�
�pt��� �� ��L�f�[O�\�*��i]���UF�O��P���_�*1�[^��h��%г_؁�fX`����v�t��4�#�J���[-G�I��!Gѐ�\t>.�2QQD��Ĥ}B�[��K@��N��B_���d�`�v�Ad^��+%	�I��F�	{�=Q_j�} �ZJP��,Ҩ��	������g�SX�I�.���)��h4#�}f�e��������l`[��1�Z/+N�#nѷ�k}{} l��-mI)�R�A�Z^_k��Y�����v_i�`�����`���(�,ON[��R�Ԁ9���gV�	ߩ�,c0K�����D�x�k똔�	@�'_���z�8����Q�1�n�n��]���ݹ��L���'ZQ!bS`H�;&OCX��l�w��*eq�2@��)H!c�:Sy��9��~10�a�`hfr���2Y�婥�%��q�(�%!QAk1�h�t퉓l|�o5*�8R�-!YG�&��_�(u� �ŏ�ג����v�� W��&=�H�%�����0�W-Q'B,;Noar�w�i~9 8���K�%���,�ø�c�^����S���z��.��!.�f�p���~�yr	�����`vܕ���5���+P` 0��&L��.�Z ����8��:���/��pH�'���������b�G���N���
,(W�$*�S��.�]���_�'Y[�Q���f�P(�i�@C_�es�}�/xӗ~�����q듒-E���������CR8�2x����}��0���_�'�d);��Z�~� 0��aR�.�����#iY�K~��_h%�\�`�D%nH5�'��`:-��wkR�_KFU�e���;>{������*�\�o10`V��(�^j��AԾh�ԚG��f���Ky�#�:��K�C�'6��J<�L,�oy:�ÄR�Z��N�`��H�0)Z�8�`֡&��xf��)�uo����\��B!�]��b颈v�e�"��2�J�aW��p�s�� ,����,��o�gn �AOԱg.%��bTX�]h�Y��;%`�B��+�h�vE]� ����;����2H��D���X�]\,�¦;!��P���Q�i�`݅T��'���0R@һ�c&T��@�k@���S�1��� C�d)��q���1��u6� �\E65@��DL�f)�,9]vY�G}��6 T]h�Nm�n�Fg8n�� ��b�^GUaA�؆r��	M��M�4�KE@�5JMm0tf+�ܜAp �A9,e-wVI��xE��m��}�V`��v�Z?b��ѼkI1�<���>J<�*u"7)}Y9	���+Y�j�h�Ā%�cP8���(���dd�,A����+K�*����$$b� ѝ]�%�d�;/
(g������	S�ޚ���� a�nY$"'�@ܪe�Ā�f-�;TH!K�niW�
SPh�j�_���t�1��v�ޛ#9�^�tMb{c�-y�z�W>�'��8���W����>/�)V`�N^�����&�R0(�&@{�D�b��]�q*蓹n�K��/_x�	k']i��e&V��	�M�|}�1�����Ӆ�Ƴod$p_��h�>�~X�� ��qu7!�u�����o�W�|��)�|��$�`K� �����;HU�Z$K<NwuH0��^��_��/���J��/��X������ ��O��)�?A'9����3w�Y7 �
��"Z���z��YN� ��)����(��	aO�bC�_��:�1Ä�����3��4+��f8��
۾��S`����=��1i��_�؃o��'�glI(�,�	�F��R4'��B����ud7�x��n���};SD���J,�.�W�
�`��M}%h�5B��`�W�8�hIpJK���鞹�M!�r,�b���Tω��!S頤:P*�K�E�L�	���b+ss-�����D�I{���@$ME{�+}�KAPp���|��V6>	G(^l,w�
h�1���I-Z��}pg�Y�I�I*�J*-�(Q�e�BYh;�^��PQ�3�i�3�/9bU��Q� WhH/�A�Z�c �8|�0���m�.��>@@�%-vX)��餠���ɝ��U iaf!/�:A�;��>�7^v�N�+q?�5[$ࢬ�-��B�!)�h	�ux���v�L���2O���a�+��g�Z�OA	�c	��6���������.�%��Y�^qE���WQh�,0A�����^2ք��hS\�>�F0��B�.�S�	�5Js����Z����\������`���n��JQ����*�8�CS�!�	��QmHgB��RhN6k�EO�iwC�zZR�%	�ٰ=(���%t0I�,c�4M�gRa<6�dI�/��P�
�t���l�1�^S������?�2�WUR��w�J�X*J��q�Y���|WK-�dX�mb���Z��ɏ|\gb uU�p��[4��r�h��	':��W~P�[�¸�N@��wO!�x��TKL���AU��SP�h�f�O��E�u		 p�U04&\�Q�����}�uD����	�7��(�.It�µ����tJ�L�+�)��6yɓd"CTW|����'h���7�V�X��B���2�U����U/���v܂`q�&/���l0w�,_sb �*�y饞t%���W��S�u֬�ρOG/02��5%#���J�R���U�<Ab&)�h8� ���_l|�feE,��՟ ��K9)��	�����X߶Y��ƻ��Ӹ�.�mH�ŧ h#mv_`G�jO�e��I MV5�=�-	gՄ�}M����VOP���w�>�)�.�ꇖ�-�K�~�gQ��Z�HP�HR�sAՃ!���~ֲ�|�w�Y�B�R���Q�/�u��Y���;(���3�p嘝p����]��������op�G ��N������ŕ�x1x;O��2��ٲ����^t��d���WG�����'-�r�`\-��hfc)���z>�/_nx��������Sn�U���Q��L�n�gF���N��'.��*'�{o�4R�[���H�%��R�y&B pmr��Z�f)�Y�Zv�^�	��+?����]R�,���(�Z=t������	��pq��ZB����o}��vh�No�_Q��v]��Dd\Z10��޴nq���C�K�J/[�1J��yR��A7g+��J��pf�
f�&��.aZh<�� ��c��;��i�¤��ۉp��pU��4e5��(���b���Uh�}o��8� nz����LL�x9��u@>��-��M/1�9(Z��>�#.1�	�X�p� �U�Iw� �t(�Q���8+�@a���\:�6��>�e%����(�k������I�΃��X�i��(h�C�L&�,���-��: Z�������9����j}�j��N��T֬)����(Te[��.����hrQz�kL�����3�y>���]-�Z�%Q]\����{� �������R�Tj`�BD`�)��o.-�/�0�%)LQ��V-�;����7BE��N>s��-�Zp	w1pؖ-�E��E��̪Ǿ�ԋ��h/�eF�N�S��W���a�� d��S�>���0�Z��L	�nЙ�aY7j���	ƽz6H[E���1��v|���-�X9Y;mv���W�6���\	��hX�Ov,��
%S^Y��ܰ���"sbP?a��k�h��K�P�	j.H t N�ց��T���w+%�WŒM�DV|c��d� @Xo+zA���U�,�pl�`���N���1�9l-����wh_܏� %�qW���P�YR� g3)�Z�� ��TnZ-���(���ʳ������q���@� 'ɺ|k^�M���|^�(W�AL����-ց�I;�o:Y�t��x��/�F# ���;�*I��bZ)Oh;>2�:p�~S�B�of��[� �~b\u�q�A��#�n[)���ۮ���g��@���T�;��,Q�F�lx-g7F�	nbf z39,��E0�X��J���\�OX%]`)CG��@��>�o�Ns7uV�]1(Z`�������u�n�Qe��JK5tA����@]Q��hq���1�Y����L�q��tF10����w%�u���lj���&\,`�Y�eN B@&9^���K�2���m����$m���.(���z�?@��`�lK��´Suͫ�U�'d�Z쯒� �_Q�	��xX}馪2��Ԁ�@"Z-�W�o�1��0��u	s|�T8�aP��	�3�8}p�	�J� G�[%[P���Tx���ĉ	��}�13�0~2��&��=��'�B�W��?�W�y-�[hH_.�������_0��Z��$΢x��Uٗ/�,d��	��o��%�-Km�w�-�t�����_�PC�ɸ�@{u9��ĕ8��b	�l�x�%�1���zŲ���%�e+�A��b� �A�M��ZD��<�AP�ᇕ��~G>!w ���w,,�hhGS�}�gN��t���[i�^���I�U+� �h� �uI2����_F�/��h8��W�鰉Jj�i�
���=��W])��4'�}�E�L��$-6@ZJ�h�g�gUBF| dtQ���%iR����N�)���I�W��TA�t:���h�J70�E#�Xn(� ����XE�OP�� ��l�f�[5{�m�����,���X�KlY�/ȑ�9)t��?�M�䞇��P�s�z�D􁯌f1���c��h�.�WV_^�����)��@	zN7���<=A�Aw4��=�&=���[-�
0��շi��2�Q�;���B���r�R�)�ߗ��:�S�y�oCh�D�@?���k���}Y_7�*�;Z
(��
!���h9���^�K���h�L+]�s�q��\s[��N1�֋���L�S��h[��gGySJ���X���8���P� h4Z=X%�}c:�iJ��'�%ؾy�Ry��S�dT�?	�������f��"������̰&�^g�DhE��>%�����fJ
�C�Һ������T��cK����������+�@j)��9O�ĸ\_OT��q��$1� ��4�z/wV�[kb��[&*�uT,���j��Z�G�:sa/�a-@�4.������ծ�%�  g��@��` u9UØ���^X�l����j�H���ך��)��KZX��jk�WG&�B�Sh�h��z�'&�yR�����X��m�,�`[E
V���L?kR�N�QԈ �ڥwb��Q�P��]�|�P\�^��$�4�dZ@��Wj|á���D� (c���2[��,�� ZXhvZc,& W}l�h_T2��5>��A!�px7������nb��w���҅�hBE�az�c�I�m�ew)�H%	_E�G�h��7(�P�ȏw����+n��R�c'���VhF\�bx� ��)�'��VDhT���?@�|�C���񕃊V����%�q�,��h�����Β���qF�/�Up�F��w�Ε۟f��F.�UO�2\����L	�ݓ�B�-{G��[���:���gM�����K��(TZUh{J00-P\x[ݲ�����_��X�@��b� ��Ғ)�A��v�_.�[�@��?}	~h�f ��]���0(�x�u�gW�G#?H^��Yz��{>/5����W�	%�A�0�JF�tmN�{��_#Dj�I��0oH'�AtrM�v�@��7�����< I䰅��]�9Z+���:O��p
2h�O@���9`H�k����0�{�q=��S��l�@�,[��	Ѭf�*��y�I6�O���%�19:�����e:h�(��ް&?G�#��+��?��Hv����@�_�7ɈQ3�*/GfY�����?��$6/�i��Rq��4W:�a;P�ŵ��b~��yT������B�X���}paA�T$�sP��L*I�D�����w�-3];�)n+�-� Nk�Li���R:�ˉ\�z9(H��Q�r�Y��}~� /�et%@�gT�X>���%A5l�~�B��=X#)('�[*�-gk��~Z`�<q\�<|�(�a^�h~6@)H�' ��K'�� ��t��e|���^>��B�Rh)�"Q���)�^�� h�'6鐟�ENT����nWR�`�/��I^��	-`\�фk���]o�lK���;��-�.�`�s0dt����馨����P�埤*���wz} ��N\�j1�j�"����Ց� (�Z"���!AK���>�֮�|�(
/�M�N/ՖK�HD[�^���,�&D��>]����4+��O�#XW��<�`�$��f��p�vдKa�FoN�/uE0M'���a�:e�oXD8JK�a��!nFڗ7b���,@x�\���N����<�f�I$���O�\λ��K����>�Ҥ�����Bk�g-�\LP>i <
S%z]gLO��L�3v�1~H��ߌ�uw�N�ھkF\lH0g�n�����0Z�f4�fǢF-��#>v�
h�+�js�B��D�iW��� )����XJe?_S����N����z0�[�V��Y�b��2_�W�X��I=�^"_K�[ ƃtw$��%Y�������W�*���^�A�Y�3/��f�).��!�b A ��Uq	f������2`	@�7���/]=ױ�� �@H� L1�K������;?��e����T�PA��y����1��g�,@�̽ؼ-PB�[c�_|���q�7�����Q����@p�e)A����$^-��s4�����q��z1PFIn�G@��[�H3��N���?*D�Ɨ�w���:� 5�JN	��@W]��Yh`�����ߛQ%�t�$.G��eM�A-��:�
���o�|K��X{�dˮ�����`�A^�0����-�Oo�b�� _RVZ���Mc��wIi�*��)$�Y>�\��ӯ���r����e7]�0�����	�F��/$������	8B�8��GĀ����\�@��W�	|:�>�yo�k�Po�A}�P|$5&���	c"�?�m�FP��cHQl'�HX<#^�Z�t(��!�D;~����Y[��� �	+;�:(�h)W��9HX<bPA���Y8S��z�� >��Ff*�%lw�{^�7�;_�\R�nGn���x+�,���d~��F�]0J�:s�J��� ��([4L����z
.3���
	���HʪBX�!�����F��^���Ԩ �N_��n�zI��X��/ 8 񥘱'�dyb�ۂB�U���-��՚�P���Yp�~ܠ�K@���ZU�X�Mz,�42K �u|
x�oUU�o�����ұA9��V���	�#-�B[�h6{�XOY�^���1B 8H�q�p@�	<�?�Z�����`��Io.m5�n�9�XQ���7��l�'��i��ĉɏha>�Y�yk��M�h�N��$v�`h�ރ�jR�	�b��z��UB�hwk�H�5��ʕA-R�:V�OZ3wj;���v&`��z�;AS�uw��4	]���$kAJ��;�vE�Ӯ	�Fw�l�&�}�U�t�h'pF�����w��ܧ�1�k�ZLT$z�O;�S&��oGIN�X�(��-�7�B��HE&O���k0v	���a;B�	����-�%[S�p� d���}
?�~�Wh�+�F�)d_�����f��́��y�ZP���ZZ�rS�%	�����F��^֮Aw�R��Hr+a��;7?1P�����ُ���.�U��j�� ���	!�M�'TXP8�jK�6�'� �(	�W:hp��$������?��^�D[��8��E��]� ��T����y�HH��L���□=/����_n��n�1�ݭi:Z���!8��c|M��/���[������h��s��3j?�D���jK�e<�Z�%����x��͟4��-�_# �2���Z�	:}�X�\��<j���2�{
�|�ǥWj��B��Y���6p8`^�a�@�Pq`"L��+�vT�)�6�ғ�{��X���X�e��Qc���V��4�7L�%�ٌ9�O+')�d�~��t��<��8�@�(����׽H�b��H�JN�-�\�v.���lD(z!$�V�FM��:/�1�K[?�	H].�`���VaPo�3RxF�i3����j��.!4:4�#�M"[A1��U�l����� ��t�V]���'�.��Zry}{�QTY�@����������/\\z0�LG�y=�)�%��`��_h/��G�'h�ir�{����ՙ.x�т��g�d`Q�9�;)J��/������:�A%��vQ�s�kփZ�1�ꧤ��q��n�>�$��ŕ�%���1��Ph1FcXz���չ�R�R+��8�O�����H�#�:i�a)�4 Y�hqͅ��	]S� �6΁�	_XKvV����B�q��H��Ya_hgn�PFz��䝀\noP�c�S���\ �C�uYh�d`��ɽ|*C�u���a�R��J��h�,�Q� P'3<�Ƽ��{��_�_�� ]�2�)-�c�f��D�2���ܸ�9A��|��;�W��K�I_�Aݍ�T�.[r�@�������iU\�O�1���Zn@�=f<�)���{@Y1��=�@���qp�re�Y� �[����r��|�%�>:&1/^��"�b�H��gU�����W���G�d���	�7 �ͤ�P�O��=�z��-��>)�^����^ݣ�e�1��$�OZ�9�\�YNU0���-H�v��']vp�i݂I1~�bav��vBΩ��K�@J=��K��-vZ`�e�%TN2/�iE���&����t�� ��@��ͰzF|��+�>~��g���z��.e�a���1�k����XQ�J�),!�J��⧘VV�$�f}bUTA[ɉU)L�2��bv_筤��\�Ta�ۓ�°����Ɛ?k��HPA.��m��X99i@��bs7P2�@�!�x�/�9U�4��t��8�m�	�]�M�f_�`�w2)��)�m�~i^�B�� ht}�No�� ��x�|�����> �[�����T���`�y��� Pe+4	� ��N�!�)�/���{1��&2�����T�䈸I/\%����.⬛h�Sh"&��p�w��H�8 �=4$LHHRLJ�j��~�T� �(��� �a��e#H��-��	��(!��Zz��_�%��F���U�Wh�	�H��gH�'L���M/����{}0�h\9:�^W�|���xR��	F�%���?���ź�h��X+����\I��'|��o��=�L�gV��� �O��'\��$FZ�h�M���w�w.���<�����ǽo�Q���,r(�zRJ� q+2>�-|�JA~�:�ּ�i���_kt�����o@L@�}�(�q �Vu8����[=9�-ʽ�b@0����I�9��𪙘/�9�>�HO*�m��p��Q�oM�qo��U%hKWF �(�jV��o$�{�,i	�l��j�K��f���sK�L�ZZ�P9�A]���2�(]_S�B��`ZhD��|k�$�uQ_����J��DV���{j ��tNJ�2K8��M�yX���xÀ�m7i�J�\v���Kʫ�gmԖ��qR�gT�yY-��z�����Q��c�#���w���b�f��U�����ׇXbfY�Q']�u���n���S�Yq�ͦ��'~UJL�&B�&u5p0 ��	��~��x���5��5�t-��o��n��F�^���'��)m�0�!@r?\��N���[Ld�^��B��{�%���`*v8yd]�FJ a�>�:��7�-�Z���̪]���|%����>BT_��i')�*����On�{� ���lOH�|��9�0�&->�'a�wMQ\@5�H��bHSt=�$��b֢��*8���7P~����~s��U�G�l��
�Lh/HFi��^+�qo��F�����ǒ����-0U
�-,��~��H�_n�1^�w;�c>�?��K��<w���Tغ��0�h���-Bn�!�1��{�`��,XsE	�y|��2	z� �0� -�-����p�e�W���\XP��E�W����Ib#'�]i-o^m��"z�3�8����~���@�y��D�(����X���������-'|Z���U�\UƓ�Z�}����Ҩ���^v R�������Ʃ�)��1UQ(��³�>��{��/.�]��ƫ7�-�"(�/	3ז��_��_V�Y��=�wE����~�G7f�U�)���h<W ���mP|�k�oO3��A��Z�K����ܒ¯ΛLք�'S�e�$���"�=B��	`|@%�����~�򴹙��НA�+�����2U�A-�����2�u�U���߫4"W��y�!�k�0�!�h�%��a�~���h�)� ��z:���@o^)�h&\����!��)*�g LC���%c6�Aj�`��:i�ب�Zbf�_HN�$T�	�H�`=�5�X?'��S%!�S�'@Iu��T$�h(٣��@�SJ`|o����@UQh�&���ߏ��q�R��~p�*c��yL<rVdF^���ZDqT+���t�LI#`|k�;�g��h^�؁G0�B�s�z�cT|���	�OB�A��ol�px-6]("���ysO*������`V{�z-=	Шnل�}��	~�R�^h{�Q�W�n�h�
�DWX�'��'�^l���[uH�w^���M�4��(c�d�Q��,�/�ZYwG��lV��h��aM{hg�K��˜��O��Rzd����=��P�7[��3�W�;F]K���X�4�r���4�p.�e
%PM����}C���P��?��]*ɞ�҉Jn�Q��,���n^�vt�	J4�(��^������(�^� C*��od���������J�`$]��iz�7z�?��5')��%��Rl٦:鏐�m/N���Y�+����{C=o^����|[]֬>	��]��'w{����h�;<s�Dd)��h�L���-�f�⢀:������R<,�,���č�'����Ӳ3��5�2�@��,P��θJ�陲u�d�{S`�H&%�AzF�|��cP40HFő��$��i�q�#e�1l%E@���*X��5 �j �BZ(����穒И���ϠY�~�I��`�0M=�z�����%W�Q��7����C��+�-`b�e��T� -90�@(5'u��J��f�}&���P�ӿ���p->��)';3P�)�ш�BR"�w�����<Y1��p�eB��_�R��k	�K[���0�ޭeJ�a{�.��\�E���	h[��xr3�iD����k��V?��b�]'>'_����5�U!Q0.�SZQ���>�hm-�.�,����m���fW��K=�	��Sl���ω�n�1�Z�hbi �l� �AXShI [-5. (�����^��]HA\�+�?FWh1,{_`Y�}"h��m�`_=I%����ӗU�6�+��b��fU_�w�>�8��>�'�-G.�.���������h\V���n�d^���{Ԗ�H�Bg����am��^ܽ}�^��R�π��i�BGw�Y0�!������< ��)�]��Mi�Qsh-f\�G���*�Fx ��f5�V�G9��`��:�d�qO�%���HM� 5����.�y�W�!R���`��Mz��7x �,-
�>�y~04.7%��ʁ�H`+�o3G7�WE�r�}��]^!?	�Q(OM;�^	��W�O2[ӊ��ZVRt^-��\�	��9>�)i� L�o����� �|C+T�r�	kZfr����S��<t���V���Q�^�PN��Na�� 6�e��_ʘh8O�����ٳ���'�t�!�?{!D5R	�|��1��siE�0LO�x�v��$$JR�,V	8��{�c��)f�o4y���u�gXQCU��P��H<��E�/B�hXT�b�&����!��U����V��]J�_{�� �:%�l	T_Ep�QRE����mP]QUh�1'�~�5���� S����R�0�ʶ��C��Q�5.��.}�����m���K��wԶ�]x���hN��_֨Q�:�z!:��m��	�~r�� ��>2n�Z��R,6�r���I Di[���`��������� 0�[J(�f���F\��[P���-�.�w@ó2�Of��4!�/�`WY�,�0�@�ag{oY��^��A�O1`Pb�i����Q��P�Z��Ke�[j�{�\h�;Q�f]n<d� ��>�Ĉk<�a�]p�_�	�1�V���H�/�א3}�k�����KnЯ�:�_L��	Q����}T�>���9(�c��(�$�~`�T��@�-�V}%�w%U� }Dh�0�� �/T1Y����)ʇ���Ta�f(Z���:�A �tPx�qA��(���STC��'@Eq	FO���d�޳EW�nH7���Y(X^8x�*۴�JB��o�[X7�;�(���>t�O��,�_&�%��镐�̹�A"Gv�j��0�ou�_ ���3�;��z���U@�3	c� 1Z��02s�uQ%��a	4=� 0"r����L�� ���,�xj<����g�6�^�Á����@ Eհ��Ee^�Ʈ��Z��z]�	�B�F��L��@�]&fbG��վ�	��qUY����T��C�m�@��Y�2>>���túӯ�[D�	%���>�*�D�@�T dX/YI��zJ-F�����]f��r�ǝ�����L��^��*u�.2�*�j�Q��,����բvP.PS�|)l�<���*(� ��T�N%V =G5�:,K�O
W��1)��Ǧr[&�<�InH�RH��zP}.J�����1��e��)�L  
�h{�a;q(H�i^3>�D���|@Vh�x�U/��{�N�PVa4�A��-�Gz�W0��(n#��hS ~ve'�$��=�&^[�7˛��Y�G8���\}�+Si� �����d ��"]I܋;�}��V�XhFXU$�;�ċ鍒W�{{ ��D_X�/�#%O�� �����ܬ]��A�k�4~����W�U6t!P������$7f��NS����"-r�H��x���'����Z�&��{�L�K0I ���`�a{)���Z������� Q�F0ĳ�h)U�9�B�TVk�#-����8{u!`h ��2XE)�W��x[+�\o˗q"�Xb��S*��sR?�u��?O��Ho��̴�
Rh�1R7As�8�@�_Keݐ��ݐ"h�g2&S}R�Z�(WR�OWS�=��Y�p�hi��R��?�%W�XH �����wX�/����n�؟��)K�'tf�]hXdqi [�r.s��K�2��n�D�� ��E�P�C��B_7'�����PE�@��`#tCxR��	y4m~U��/�7�NX��X-R�`}��W�TDv�Vt�м�$+`)�@:S��~�����_�)��82�A��"��f"�H� ]�w�D�|`�)�/�z�f���@[��/���[�>XN^�JDQ��Ҩ#L)wԒ"
O^�Y�� �i�\������0V!p(�bbL�F�Yh��g7�Х�h_Fau�N%�B�ݼ%V�R@��"(n�%�Γ���ȣ�=1G�Mҁx-�c�m/�&Q(hr�)�����TM�\e:7� ?h�E�1&Ո��{�	�H	��G�|��j@'h%7i���	Ch�^�a5B��)+�^�h�ީ`spu~���y���9q����g��䭞��t� ��hY�յ�N�j0|`g^K%.�U��%�)��� SUh}']�	9%�{N�0�T@�Z[C�ڸ
	�D'
�L�- )_	�(x@��A0|mo�c1X��"ijO�R!�Z���5L�/���?Ф�V�>Z�7g}���j^�����K��� <�l���(���@�=�Q\�J��E"#.a5ӓ
d����J���X:�;�2R�)Y|;ky_�~���<d�	�'Fh�����-�J��Xʐ7��uI��h����!F#N �[�n���H�t�&�j/6�#�4*-}��d�!�������bA���W�0�U��o���*f/)\�S[��B����H|������������U�x,1��h��k�|/@SZ�~�RA�+(�Pҁ����K���QV�(���aUy��$�Y��`*�C��G�h��' �FG�<Q�7|o%^	�D	AL ��Q�a�W�4��83J�,l�Zl;	���H�r�}�^�퇘��g,�?�% v�Aa%�-"�L+6QH�?���	H�Z`�\�d ��G�=2 ��z%f���NHD".	�/W����W�Zq�?&��U�2��i��੸�,�\��]~��(X1dk G�e�V��3�;&-�:(x���{zA�D)�	���p�t�{����
F�<D�\OC�MƲ����PG��S�������5��5LWFrWֶTv���B����V��,��&�� ��1�-�^�I������XR�%�Q�it͏kMa[��	?ڮ^��r{M�O�h�[h�o��9ˌٜe .dE-��1 @HL[�C%<^��ܹ ���7.g)�КH{ k�&��5���~�nwI�t	nL2]WH�l'�{@Ai��P�d�)��0H$�aq �lj�K�[֨1��_�w{����]-FKV8�����_��\fq��2���	��V*g���-,}��-蒥4��݈�X��nZ0�fKHRWoү�����Y�o^�WPH�I���L%׺ ���.RM_=�f�g���A^~ p5L S��N�()�[[��h9. ��@Y����ؼ�-Ѡ0��|���Q��#`CU�O	}��X��A�~���fXWh>S��5Rf�%�A�S�8	�2��%_B�+�AQ ڵ$I�|] T_��п���zU9[�� �]���{���00�x�I�w��K�dc�����- ���n��}QhRL' )�?(�L�,�<e��&[ZS��7�vm	�
	�r ����9��V@���/e�]rO��5� ]S�OM�~<�K�YK�fA�.�rz�)�^�^��V7.�Eg��k���V����(�stc	b��1�ɝWo)~(�;@(�>�͠���%��P�%*bq��cj~�#�x߰�A�j��SVc9/Y�,f���]���0_�V& S@�n\w���W��L�-���e.��-�	�Z0g�N)���8�н�9�t�z��VXZJ�s���� �-�n/X_�9N�|/�[�*�-hf!����8�^�X<�醚�?�K,a-���o ~h��Wa}3tc,p�|��hMK��$���9�`����Z(��ƫX_�U��=�I-��`Q�3�Z��/��g���� �Hd�-1�_����P��?�[� �¢�L!X�H/ H�^@9�Y��Ik��q��� k]���xH���e��[��@(�Ї���b<�F^��؁l���7.��k�@��6���`��[(�Y�����G�@S���w�:�ˏ�RB�� ��%��jfho?��d�9/S+��#Pp ^O���G���^�*ř�����.��,��	��� ��YM9[*�
��h%dff�%xDc����P�ė�G��wA�(�]�C)�DT,
YLI�'}�^ZhH/�_
�/]�()�� ��K1n�3uPtV��$�E��n0��"%q@x~�9t�%�L�O��ۉ�']G�R*���;��9-\v�r�>���b�&��s�K�V-�VHZ�ĭ�[!���JnV��,>�:qv|@�<z.�#�!�l	�m�/�d{1�&[��������w.�*J��e�
gW���o��?�6vO*��.�f]rʑ�e˄��&Aj(i0_vZ�<���Af�J��8�)@�1� 52 �X����A���^V��H^���K �1e���Hu%	Wl�-0��[�����9�>����Լ�Iwր�+a��?D�Mƥ�[<��%���)։{�(��^HJ>-��'�Ku�� 9� ���$;�G��:�`�����k�1���t`���D=dg����	N�=�;�[��@ܸ!.eU��;G�>�%�v��Z�X�	�K�$P2��^@�A�Q�,�1�L��
E�׉ք�K_C30DL��XwyQ���9�r|�iw���x�!��B�[=�e3=Y#(�,IT%}����,�)�.-HS	%�c���n��ܺ1�(�Y�2A1+D,�S�1+3T��z�TR��L����	D2Ja�y߼��fv,e3(ˣ��V����5D���礔G�+�o�y|����XŸ2�d� ��F1:�N[^��w��m�v�2,�1
QU�o��{�� E'f��p��R0��N@�^^1�B��a���W�즸�Y\���0"��S&�Hj �P��,|�j��;� �҉�7	^k"E_�?Z�-$��ʞP�S;�T�ږ/8�ŗ��yU`�R@�w�0�<��nH>�r��(�NZ�d9�(�f���3��H�ƿI��0/$+�#gAB*�5=�K�S
b�'��x�cv ���V�^�w�����8 J�X���&\^[��q#�}C(�a�)`w�%sz��Q%�),i#cUB�Ut�H�R�::#�cѵ��sߝJ�}bi��Wb�+�- �Y��h
������E1 �UTκ%[ռ�%�!<{�`,gk�BW ����
��M*hpK�UYd@&�=�R��N�z�]��L˾0�W�.��'�U%X��}YZ���)7ے	�i��߻#Q��/p��3�]�V&�0�b���Z	��DL}���R���	��6��ü|Z�u�hhڸ�U�񄃺H�o��,ܥ1�H��V��(�B���ٓ����JH'9��A0<�@�J��^B؂�KM���@8�,�_d��a�k0uh!�aQ|�>G�ϱX�N�hsǛץ�)��`	�e����^T�]-�	D-u�%8�[�)?n�a���+���)�l��h>'n��N;@1�ߚ5w��h;�U���Z�=�c���RP����X�Ԡ�yH�)ט~u=��Iϐwf�[R�o������H�����Z��zXҶ(y�k�-f��t�
����!K�"��Ѹ%$��yNCĄ�{�E�y�'h�c->Jy�%�`xv�]|�OS����V�]Z���lOmT�mZ�V@C�g' H~<Y��i��'P]|:���(�Ըx�_�"��+�����v�H)���a.��C�-W��ґ�;��5w�� h��3B��|	��]3	[4	�������b8�� 2)�d��x��H�1�o�:�tҺ�F. S�ʀ���;�sL��N��@"�J
�h���Zǈ�J��S�h�NZ�2|�L��hq��e���ˏ�9TB>��G"�H�������ֻA���1;4CV��@�]O�O���P@��l'������W����0�<��Ubi���{A�U�2�7��u<<,���F�{�'r����?fh�﮿�a��?w�RysfSL� �ہ������+b#b�L_�5()���S����%��.�PhgN̳R(v~��Km��Nx����b��7d�?����OY��(_�����K����$�>�z�e�b^�MO-6.�,nVF{K|�	P~؝_\�q#�o�'�����W�\P�%��*����+�MU�殂�:�����+�<�h/�
f='��&����b ��ᆙ'5��q(_��yR#��C>
6<�̀� w[�m��^(�k��]gX�R�,-�r߀�P�qk&�d$$�����}�y�c����vA���J� *�m�.�;��i!0�Yt1�-	���<�z�
O(�5L�x*-���x b��;��?�FJ_���2�qW���,gB����,YA��ĝ!���l]�?�+g��{�h�w%��|/���P4��kX5�����u.�1���
�$���:��Vc����7�M|�a(���_*��� q6)VW��%L����=�{F�r�&��m�޳�#�cN.�P5Y�4���6�aRP��0���\[8�B�\HۺK/PAg#Q�z�K�R_-���GU�7��8����oRu�R�h{����r���4X���E�	�OV�o�쀓/���V̹����7�͇Q>��2	�:��
OI����V��F(��}�7��ј��lVh�.<YdQT�8��p�
RX�����e��
�a&^G�aӹtZb�]X@� �%�K�k-tF�&����_��K�6'
K�X��'p�\`��^	���jq�@�fX�M��:|��<�� �)�����4r�mA��nrR�.`Cvנ���L�5%D�<��h�5�e�U���'�܆�Ͷ��a�* �)�Y1��_B-;7�J�p���J4	�/�D���&M?��O��;���/z� =JI7J1�ף:��?�QyN�Vv���J �j1�%�U|ti}Ե�^M�e�(G�K��Ҟ�ݰ{�,Z�����)F��*��Nj�J��;W�j�t�^������[��ǹ�c��+�8V�F����́��y�'1͓$��lj�@��)�#��X��ZV�Z�� Wh~b�T_�`T{M�a��2gBt�	#Hn�쨚C�K	��ҝ�W�k�v�-�U��`u/<|�� ��D���%�_2k���(�_�X�yN�%��)��
x�tV�8Q+���Ʉv�[���7� ��Q�{m%e5���'���Owј�\�ؽ<�~���r\�4�xXW���	�_S����v�%���YSV	>?)�j��ϔ��1���P�� ��\�-i�uF]h�{�<k�	����`�#.xƧ��N� E����;d�ʝi�X��ǡ���A�h;��^�D�p۪��"���'� 3 -�>uT|FW�H5[���))��,�EW����0*C�[Ss_M^n!v��U ��q��e
��<1�(zV��!�9�r%�^�݋7T15��X����%$[�A4{��h*�IKa�鎧>��T�=U 2l}�:;�TRX%w<%n����,E�	�/�tiT+0��'��u��^���L6A�)~�%E�L����o,WEZ�cr�������u�B�d�%���h$O|�o�H���҄��([s����/�GIP���?%{�f�r��L�1���h��/P�����f��h���m���6)�N��-	��S��h�%�WıP�CN����_�.�R��>&	�)��ThiO�4f� ��	H,P��Y:�2��x��ash@.A:��kU��^��,�C"��;�Ŀz�����E��2�6��Cer���Pl�}%��Ĉ��
E�T0.��}�$��B\4�lqi���Q˲Z��<�� �����4!�u���r��P��2B�a��<����Z$^�*����*I��}TC�9@zCu����i�-Y�����;+�8uONR7�:��@���O|�W��a�m] ��t=Fc�dѰ_	y,A�X�
�]����(?	y�!���5h<Ը5�2��BR� 4�9��g��u[E�U�q�l�4��� �J��!W@�4$ug+e/��ؖ����V%R�	�0_:��X����	U����Vm�P0�X]U�h-;�)��}_��-J�9��s	l(4�(�,`��]/���`��I�X����aj@n�\�!������넒�qeac�����ޟ��_�I��%fv;b~�M�K �U��>�t���
1\e�7�o`��Cb�s�c+�Cӫ���!��
'���cR']w� �.�"HS� z',�~z_�XQ-.�Sh��3�bl�/)ѫdP�/��J�}ц`�Ԁ����DV�@��)#s�O͋�N��O�$�{�U��B+��^��,�[�+ ��-�)�8�F�}��DD�T�j��_܀����=p�w3���*�Pm���{�1)�E^�Vz�v�E�B7� �S���� �[����C��fSRA�Wn�<ӄ����b�K��J�80.�N$��`Z@��k�=����n^���=�Ao}1~Fq�.#�f{y��Z)�!��.�lI�X7��)=LoJB�i�H/�5�V�4�v����Rr�_u�WPF-=�y���	��ha\��-�DI��ܢ��� ]2{Xh%_�m���(�4k�
8�`�������0���m�+�o��.�	J����2�X>V�&f+�T�������Q�X�j�i��0phM��a�L��LL�������^��,��f)}
@�b�	o�1�
3���b�T]�D\����q���	�V����AU'?r��-�$>��{�E�	IVs%���A��^	Kgs��h�c�Ե��P��\{��rK�A�?k):ڱ�Xn�:������A��d��I|V[ ~���� ��^ބ}��P���:�7�U6>ټ��/ER����^'	�zwq�o �^a/��Z�Q-n؆�Zl�*�KD�j` �o8v�q�	�eN@�ٕ��DN���e0]1�AB�9l�/�L-��%�V�t���S��b")�UN���6STJ�a�>=��ɕ;�\px��4�	G���/]���|��輎�Q��1= ������sW�y���s�=��q�rzN IA����时TZ�x�F����fh���t�USɯ��o��:�e~X ��(F��C�A�l���Y�i�J�˂ae�k��������#(�Z��p�L�7[-�٦t5N�0~I=E�w�����?�`t���K��QO�A�|���c.x4:I�u*҅�ׯR_W�A�F�4넌��=]°V�7.@�	J2� �%\/��.�TJ����π�WhnNC�k d�e�x/�R�<�,���}�n��)vy���J&0��y�E�*���]�-=n���T�-iY�ˑk&�T��Kb0*�} ��L��(h�� %[�K�4�3�z��V���O鐉ZL�!+\�j�����ͦaJ ��c5'�O~d��g�>���!H%�2�5�X	� 'o� .�G;FJ����w
^��v�_{�,��=$�/����\r�m
Q͍ڟQ�9^5�u�����M�H��%S�9!`�TC��Z�p��4� 3
��֨��D�{��
'X@N:%�.� ��R�갬����B�_#�㯆{Ϳr/��{�!���h�	�氒�!�v.A9�7���@��r��V�[B��ҌJ|�[U�|��+�b���Yvu��-�0"rY`�"~�L\M�C�v!鈸��;����aa�ɧ�ΐ��K<3Y�љ�����D&kH�bG/Y{	��=���� b�&����8`��DS�Hj� v��1�:���h%c/qÉ!W41_�x�)�?���R���	o����}���WN����5E ���U-�-���0���ik��}�ZaH��BT^����Ψ[��ؕw���Zר�׿��YwE 	�X�'Xx�I�_'-�����(�s֮7R`�
��8/u�Z7K^�E�j�Md5���vy �s���[
��+�R��u����$]V�O�9�h�X�l��
,�!��B>ghu��T����)��*��U1�k��(q��C�~�	aDD��n��S%_���Y�#�Ղ�]{h��p�����?���A����ݠ+�Ѥ[�S�	�@rq	�ꐖ*��z[bӜ�DI����퍧�,���-w�^��~��	��
Z���R�ӞQ�i�^�Kb�P)D_��?����Hӫ ��*���,�(��� ��"Y`�Q�}���ǝ$!�X��@�V���9A[����2��I[��o֔\+	����,�1}�ZQ�M��%0oL�ϐ%�Xv�Rh�>���NQr\� ��@��Pi:1��}4����-�z��3l�C!���"	SP��p��HV��¼i9�î�� K�����/�<��R_Vg�鵕�,�2J1�Bpm,\� *-n�mE;6i._P̠�(O����6]���y��5�hV��r�_+��@X��ωh��f.'��	KtV�҄��R��
�u?ƻx&�%�f�U�fƎ;����)N18Ef��-��.��1,N�ldoT����Dh�I����aQX:�aL�K�Aw�C,�2╮��>�[��flڶ��u���?Q0�fZ�k��V���ҮD�?�T���\����mx��0t�G�O&�v� 2e\Z1�NXƿ�gj<�GR�U��#���'��<��Cc �摀	�^nh��ݗ���3�8V�nGz@���f{TI_Y�^)�ޔ�=�Gú����@�X�bW�۸��bS_P��'	RWsFe�q���(N�=�_��h��<�D8����-�"���	]p�;��'��� E(�R�O�e$Y�.O�(}�/ؚ���2T���hQ����8L[X!ǋW.��\P�%!��0,�7�Eڰ}h�l`D���y����m�^.�%+��B/���D%uFπ�"~3���pW4��@X��@����������o�f��.x@���\�ɀ�ŧ
��������Ձ��u�����ZP�j����*�n(�X0���t�	�_��'P�~;[���*�eK�.1 	!�h܃:� ���J ���1|�'-��������ٯcN��: ����������J�����It��nW�6�
\_��	T�p`�^?�|)��W耷��n;�p��?�lUd#��nW�
�m3�}��=��;����ac!�4#�L)'ԙ�V+a�/�j��]h�d�����+퍡�,�2Gk��e �NU!hWs������O�1J���	�����b�p#fL�Gb�ՋVV]F�&���`�4u�(�X��N�M���N��\V--�]��h�7�=�qz��0�r^I�Ž0]��a9-}>^��X�n��y���q]GT�:�a+� �JE�H<��	�p�%S���9o��-��:"L[^�?�b�]��Qfhtp e.N��)�aj�_&9�z�OUv�I�G-��Q�;���r.hdG����U�6�_v(���hX^�4m���t*���k�
�儰�������h:�	����`z-�]6�7U͡4H. �^7���J ����^ ,�X�G@�}�����B[d-T^lO��RK�PBI׀U��	*L#�9���U��\a���>g�0��2�G�����{���'q��h�F�^���������k0�m�Vh�p1��<�;EyR|�3�b�_��m�:���r0�Cxf�k����o_VՈ�:��0|�	��|c�K1P?�ϵ�ʗ��R섗��TWT'� ��X��Bm���bÜ<�]1ؘ-�����vc�_�e X-8Á:�E�,l���u��-&4�5�\iv�H

R�-�-?%{��K���rJ2=	/��P�W��q�&�%� X7�*��}���3L�0�^��'(��ȋ�5%����/�@�fe�r�@ HQ�$���h�m�2gti�Y?y�z^�lXb,���BzY���O��B&�ũ'�|���:�!��h-�a8]p�INs��&N@��%!}��0��x�����-�n¥��¹v]�-����݀�;bt� ��Ea��+֥�w|;>=�����$
���C�i����b}�]�q;����~}f��\�Ӿ��`�Q=
�ު<z����G9^���� -]�ww���{X�⛨�Ts>�|�_�>h�Ǵ��Z&k|46�|��F����8�A���C�ew��d�O����m��������b#_�g4nI�۪���	�"�A�y@)L�-%$�_rWt��U��wh?W���Іt�"���i�5H�`�L*� VPhq�=�%�	�e�r-K���i����ޝ%��0��yR/Ob���J��O�&��KX�a���������K�_��-�Vh�n$HUwB��u�5����+?
���%p�{�C�J��
x/_��KDׅ����� �O	1����^�6�QhNy7��l�,�f�Nu��;	���H�P���	̀���PDo{B�a/k3�~)ΓY박��v>����n�xq%�|�u���T��c�-���n$�여�0�.� e����M]E8�l1��]f�x'Yo�I}����D��B�A��~ڽ ��W�$t�
K��?_��J��'�Bs�qr��A����鋭�|u�ܬa{0%M��}B=���5�N���ac�n�R���e�|v���������3Ls���D��Z�NZ1-�#��M¥����՚�ގ�]Y<�wn�uK0��Hu��!���l^DF|����	�7UO��� ��Ko�k�B|~V�`O	�^.���/����J=�%�+�)w�M@q^�5o�_�@���f\��J��;��k�O@�\�Y���8�_t�P�o$�jU�3ɼ4�"Ih�Տ��ew|y>�`Si�!
^GKspNP�#�PP>@h	'1{2%ޡ/�=���h�2�+��}(�)_��)W{|��ے���Z(��⪞����h���2
~��^�1�d���`v:��A�Cʝ �m�3��?�M����V}y��Do�E�.z�š���\JFaG�P�1%�0��A���1����%N ~5�1ix#L�,j�
r��1�(a]�W�2�"K���� �w���3@�a
�j�<O��9en�ŕ8	h�E��W�I���(�iϟ�s������H�6z)J��h���f^���^���X��;�ګa+�	�|-���"����ݧJ�{/��� "H.)�H��� P�cL�?4%�Y`�>k}Q��Ӕ��`Im����ah�`�.ߓ+��,Z(�h-GC�ø�)B!_��W2&^[���?����P�~%���Ű	%�KS�vJ/�A�U0}Ja�̧�Μ�Z����P߅n��z�_�-U��:�NtW� d�����(R����~��^-����q��ϐYq9�����%����70�|)��.�\��2�QC ZwG@^����	�1��+��r���K����0.�+/NQ�ܻ�cq%��Z��3;�����첯8���ܞ��[�F� �Q㝀۴R�t��x!e��q��E R�Z/cR��2�S)T.���+,X.D(O]���)/����ŗ�!���F�-"�D��z� ��Zp;_ ��i�J�u ���z92��H\���2Udr}�g/]���3R&��wP����%W&p����[~����2���%��	2Ww���.�_G?�J�������K��P�����D��`4-�&�'_%���, <8@)]3XQ�ɥ*����W��Q�dP��\p�?��`aY�P+��$&��'���� �a=�{\Y�~����$�� &-�N��3��rӻ1ol����K�M=_�}�K��0��N��v����Ou[.��ݟ��1`��-��|C���X�-�݅G@�:���K>${�0���!/Or�X�G]�5�zh`����d���t=Q�|�5��X�%�E~pr����:�ut��\�����<��7_�b(��Ru~�ah9�_�¡D �)x^Hf�7(�߯ڶ�з�@S (�_'���o�W^��օ����X^-�e����U�!CY v��1N+ )���(7���	�'ѷ,��P������N ��NC)ڒf�n���ƙ7!�C�(ZT�	��)�b��y�(���D���8�Fj��k �N(2x�+t��i�C�~��5���7�	�q�!��V�)�R�ZN ������<L˩�K���!�M�F;⥗p�#�h�6�g@������P�ǿ�e�+��Zm�8^�wR�{�\%���X��Sh-�i�w�\�S�If�{��o����^�}O�v�QL:h�=!(������սJ���[>,�����������D�Օz��3	�]1L��;<�~O��{9��)��hj�[��S']��XY>(a���������	�{<�c�Ӻ���Q�"�W�e�78�@P�G_������QhR3�J)��J�2��H�	�@{�.0��@k[A�K��#9jr��J���,lqA1~��-�\b=��t�.�0]�gi'YPL��;~�P,�ߐ� t}L���E����!j~A=GW9;�N	�(��E����dBZ����)���:	�_r)���^PU���+�h0Ԣ_�!�;U�どYh]T�� �ot,Z!&�]�M��cز�I��z��[�x���9�@b/3���%�w��� ����0�Za����G�S�%��88@Ǹg7����~S�\���j��U�0 h�Q������W��^1��)���}6z2�P��hb+�Q*p$ R%ei�c�����/�DĒ������('R����]c'_u*�C�}ؕ,�K�O֭1�yC$R��ؽ �63��0�qz�p�)�!Mj�N�e�˹F-��/��T�� Z@M-4�f��7Z�(/�	���;�VG�ʾ�Ri�JD�2<��LO�.��v��{�ͨ=�O:���e�C- h�[��`V_%�I�����j]�;�+	}#/oI�_m`���_��X_qwk�}�.���-��j>u"��\�`e?�(U��p�'�.w���]�;P�ihAIb��)��� �	 ��*�.CD���� p$����;�~�L˰�� ��/}sf��O	)�P0�K�d� B�vF/i� T�4"k�p!���0^X�ꤴ�����$��%_�;9^3�b �YO1�v2Ix�F�����#����
=�c@	�	%W��X��<x!�u g,'��h8-������)��1�>����<�$����ci�uPذ5�-�r&�8e��ڈ_�`	�jA�J)���=�A:���{�8=�����vQ��RROYA��1π��_P	����B����h���u��h�q��髴�����3}�$�����k�[}�-��#�(V�y�T��-�~�u_����2�Ta�| ��h[E��<���N��dzR�	���Ŗ�J�cؾNή��J��O�,�@.h'�_�X��� W�1~��ןT�l' ���u��7Z�G�B+�Ät6	^�s��u��xR�������Q��(_���IT^Y�y�/]>�Ԏ�9�X�9,�$Y�	o�U�������r�"�V\ɨ>O�ĵ��iAT��-�ĸ3HƼ$��GêG�� ���o�j�A?� �h�N+1�0쁓�\=?PEZ�F�Q"�|�U|rq�-3Ln5�4�O�	\V,`'����Y�uB�l=[)ˬm{'"J�
�U-%#�ch*�3��!"�4�H	���p|(Հ�7�qZf[ofλ���o�<����� ���f�P�V/�r b`d� �0��#��l/31�_�@�.�A����	kc��������[E�����|�YbG�먁j�S����d��O������5�t�Y�樄�[S�PI�j �G�P
��.�4�.z����y.º�����kRW���"YW�2K��Z'XPn��R<��XA�W�s	�9~�ꖫ�5N��{�
Yh�J��Z��]UEc�J�T�M�d?:H�cj�'E���~��{wx@��*%)�<5�͒ �����fh{)Zs��S�Ƭ����;p@���-^���L���I�j~2\�x,��>	���2�L 3g!}�����%B��(^��\W����%
��Q'�=>s'Fr���O�D=(�Q}z���^~�/-�	�����2����dS�����鶈�%Vfi�M���:������-���֮�@X��h�>�*^������p.��-}J@�� ]%�<CH���>S?���S;I�Cd�K�@��k����h3qu`�I'+&��@�����:����g~��3}I(�鷀��Q�|~V��c��hz��f��-���*�0{�ʻ��]��8m���?�s)f2��_(��`�`:	 ��;�H1�_�v��x)�>thUeD4���_]�K�wDs����+�ʀq0�T-Ɍ�+�PX���Ry h�b|^N��i�>:`���EHy�L��ŗ
@��G^����$��|id�N)��&z��=Šj�Z�F����p%<������|�Rbi|t��*�P�omK���<%�i4GH�^�f\���f��Qh}Z�Y���J�����~u �-@�5{;�0��~�EJ@�Z/4�Cզo�	{��@X-hl�� 4r�+�֞�z`0�0���]ѭ���n�΀�!F�N&��[ K�Y�j�@TJB�h"F���1,yN�q(���*`��2$su{��)�N�RƤ͟����f�@��0�ېt�_�����	K}�%(�m�&"/�#�=\[#�)~�B�s�Yb��4H~�>j���b�fPҞ$F�)�d��A+s�'�T�b�I�y�~FXK��j��ī���:�)Ey5�����U�+�@h8/\O�i�.� ��,�`���)���̕6�� %f��-�j��l2%tؿ �,� �sxg��@)�Z_�� 5���:��w�˫Drhqs�ggA�'>��T�蔬���x���h	�F�	�	Vء��l	��t�r_���}*�h�v`���oB{��;��+Ym~�Ƙ��W��`�w�k��]y6T �]���Z�%�WAp��_	x�%�T�b�D�&�L��N�
�@3�����w h�1%Y�̲��Z�oH_@��(�[I]��a���H��.�eV�<4�,��'UF�Z��h2���%��[��wн|m1�&Ph��K�O�1�/R�Y;�U�H[?,T��;�t���1L
o�:����ؿ�/ax��~�M��`�{<��O>�L,HF�-�$QEGT���>ZY��OD^��<|ǅ�M�FK��į��Dǉ�,/F��P&֝s�5���M~���c[p0�r��|0Q h�0�Q��X���T���#���E�,H h`A��bCT��9�z�䪩��]VQVN\�������L� o(�[nt
��[`�����a^"�cYhm%_E+Bޮb(��E')�l��YLe.V�vy�7�Lv	��Z��A�Qa~�6خ�J��%6X�JY���>M��ҭ8����u�^�h�IW�Mk(����a���/7LH#?z�*0��&��)-�D�l��K2쪤�!x֨v�:;�K�} O��g�> �EW-8��1ºd��.7��+�c�@SZ�\꽭�c���_Z�9�����(�	��}�VN��QbTY`�������TG���uDPe}k౔=���gK�rJ�V�I�)h�(��>��w���R)��O�����b]��������;Ӑ�&�A�v"cw�����i����V빴�F�xf��[)�?�	���wj��׮r�]��;,���R: �8G�?�U�#��]~�BpEvX6���D�����X?����D׶0�����u��1}l2��(vX��{�8pG���̂:�G�C��V~��? rp?W����f���{I�U�:�<Sc'��_e��Gh��Q��2�Z1x�TݕZ�e �N�D��u�;��iB�����߯>�íz�
 ̻�w���}��M.�{�쒄G2�/J�����}|��%���uI`-�!]<�y�������`�Ŀ�+�8�����;]
�3��=��l���;pw8�攢���I��6B)�5{%M&OZz���N%]���W��o,��&qS|ǧ�h)Hn���١� 9��̍�C`��]%^�T" ��#Dt���!r�6)h��Y�HX��4�.�Sfx?�Y�i6�JsX�� I�U������CvR�Q��h4W�:��{wOy�S�� D)�[���>O�(Mh%�p���Ft�9���d����-�陊K�5�����[t��!�6 �f[h%_W�4/��$kO�bB��	] ���5�Xw����ܐ�n+	��)�u؈��؁�u�'�f�y)����݉CARA{5|�SH� ���=�@���sQ%��բO�j�f��3���KUHW΁W;�����SQr���?��G5�n h��y$]ET'�N�=3��^IW��'�������|�\���E=�l/��	�a�x�y�������
������x�DB�)K'��}��Z+"��U�/��~�SP9��J����zN9���)�[,��b�Wf1zxI;-^CR���L�'x�����v.��2� ��\�+����n���'騷�1����iV�JN�)Q_Y�|�$��\%�}�E�]kr����F/X)��//^�� ��E��I��	 �ڟ�u'���wY�� X\J�i6o��'� 6h�]\�:S�x*�3Qh���%1�)_1��ߘ���j]uYą�r��4�q��� RWZ_O������e�!��"i:I���#*
�����H�h��-3����p`�h�F�j��/CT:K��X飂m^TY/\=O͠?�eX�l!���p��a`2{����(��j���3��dc%�ѣ���B`^�:�i��t��d��eALo-Jp��]P�4�ZSڬ���@�I��l-Q��B^AC�P���[}�aG���O��?z�		Ok���	u�vD���n�J���PZ�@Y!բ=~�Q'���[�%Zꁠ��t� f�r����.���*}�3��:MF��y��0��k���_���%�1�D�^�;��`@C+j�l�yÖ�b[�]��.!�B˴_�ab��J��y�����HZ-�J\�%ՠf��e|��&Jx����Xq*DT���n�b��h�9$��M�XJ�0������t-B��]O�:�DA;�:<��C12��8�d��O�'�������42]�0	�aZ�c�z��*0��V'��S�-"#:�h����r ��P��y@���N�f	]Yn���SJ�- ��p�H 5Bo�b�?ڔP���"&T/�_�#p[��!h�.��zN{,�r*�����ie�vUC�K)L(�Q����+��:���^��v�R���	������%���^df��Xb	X[V1r���M+,���� Ɲ1nJ-��/��:O����DYuD�h�'�	�U���7�ya��o�F��g2MBXBY��<��ƴ�Dw��R o�g���7��21�T�%Ցv��f��V��_�p��8�!@�����T���+(������8��yM?@W�	�[�)V8��Hf��9��É �'D�O
�d�X>��A�+�d��ـdf��&ڱ���
�ؘŌV��I�h�[�h�N��R'\S s�S�GN,ȓ��K ���phW�o^�D�D�G�I*Iz�O�e����Z\���7V�����$��Z�\R��>�2�8��A�o��)�u�`6�ͼ#EO�#�ݨ��,�b��-&���.�Q�+�e����P���(��X?�����;$���RA���@���į������Prh^DK7<���n�i���3�N�㟣�[������������=�J��� [��0�ނ�݀=����(�<,}�xK�*0�-./�j�  ��{ ���i�P�qfHrZ{$y�p�+�b'��XA^������O8��Kph{�;���@�Y���1]���z������*�*w���4�{5a^o�J�Ƕ�=�� ��gq�)���|�EP��5yrH.�l�A`� 1/N+��y:Ut!�b���3#p���b���N^�d�NJU��'	�F0	�&' ;�j�Hh N��	�H�u�9_�w��(	5o,K� ��/~K��-�8���.V��i�Z�d��<�Jh!�p�N�Bpg'��Q�&�	"�s)���,8��}�,T��w< mS;_-M7|)� Z��h�[n�s�>0�pN>U~�u[�9W%v_M��t�������{�0�p���!-T��o��8{�	Ř�@�� �0�]���.�~0R�F�vu�U�<�K��\XY�ߺ��}�.[�/H��i$Qǐ!u���U��V���^�GT �;��~�Z��ai�w��i�N]�w%�1uAWY>������ү�-�rUB@�=��ņ5�^���P�m�'e�p)���E;�sΙ�U^
HԐ�'N�lN���e���d���8Wh2D��-�'W�LX�L�O�8�,���� �c:QT�EM�\z)�@���9B�hQ)�F�(�<D>�]O�0��u���Uct�lk̳@2h*_9�-B�y�Pgͩѩiwz-���M����A�gB�w�6^�q� ������d�]�����]�O�\���lEN����$�k|�&z j͞c%2f�xq �p�{�
J-�7֮���6�-UA�.>E�B���aK�]�途o�/'[�<�%f��I��@
?�}�u����^B��J*��>YU3�kT���$��S/AAho�	ai�k�tSh�tz��]��6EKi+ kQ�4�� sxL:����%�e��^�X��f-��{-)\�p(y��-1��#��{cN�铗��O��g
���)U�����D�`dR�Y�����+���hD$~�S�0Xم<*`���ǋ�faU�̐e�:gh�5l1�\X�iq� (�����,V�Yaځӄ��BK�T�>/��,��fR�3;0�Z����](���Hk���P<^��k�1*QV�0)�B �S�0��d���ػ�h�%u'v�q4<q�4�a�@�WЄ��^Z�8���Z��ܭ��ah�:&��qrF�<T���'�|s�=�8|0ϳ-�'mn_D�*����^R�'^���{*�fKPJh�)�ry�=��ŖK$�)L@��AR2k� c%6-����_]_	��O촚�Xbhr;>	�.����ԉ��_U��N�$Ʉ��OS8l0[	/�l��1�k���dI�?$:ݺ1�G��D���ªN(�%�"����Բ*���?7{�����'���"�U�/y���2�i]��A�1�^� i&w[B�_�E�=:�'�|�A��&5�L$��[�I%=Cj��]항���\�6�f�#'_t�֥֟�(����/ �e��!��'��RB{=wB�	�������J���"��� 0!�-(Sh����J��r";��y�����3�z�
��H�$TN� M	vw���&(m��U\/s{hv`��8n�d��OǗ����F�]�咀��^R�h��4}�l�m7 X���+�4\�l�	ᦓZ���^��B�F� �6USER32.dl<ADV2PI�NT�L�T
x9E���o�(h��
B��`L+���B��$�!���q䉿	1����{�H�����������a�������78R;�`< �9Q> �e=i�:L� ZF���d` �"�T�*���� ��y�.� 5J��N�� V����	�8.�8���ϰ�(��]�ܐ�!� �A�%f�� ����� #\�����8rf �x�r=k*�wK '̔���="�>�wa�^�Q����+$���y��� � *�R�w� ��b���� �����W������� �@oj���G} 6�/���� ������@E��v*�I�p��������� �8?Q<�_;Pa�R=�f>h�K�Y(G���e_pV�������d ��W��) i7[�%n�� ��ksE�M �`�i[GO��?�nǀ6����$��U:�� �6����3 w����8Lpq7[}5kr�N��\99nA'�p�3+���V�Et{OkȒhDluUmV��Ep wSڝ���u�R��������P��Ty����!���RN���<s5������&� 8[�9}�	C���J2_ gu�/���]$��%�@�1�F^D�GY+ h\��L��� ���H�� Ƶ����� �����؄��U��f�,� ]�V�R�gwh�Goz�������.;u}:�=�i�U�j ԡ!�Z�$�`b�wb�L;{9y'�~���6���,n&ç1!���G��b��p $|��%��ـ'�Ӹ+�U�,Q��+����@�h�\̴� /�Jl*j6}(�;� ���'s�M �YiU�\X?�QOw0� =rHdK�E[`t�)�`�i�`�^`B���(�!�a��v��X�l8@���+��<� �)�*����'�q�1�PͰ� .�(�[�/c=��x�5 X;�UTK�☯��w� ����C�3A_)��}0(D���	�׿/� 7cE{� Rf��)��G�s�8T� Ű��	�9�Z�D�S���C@w@��� X����d ��	�3�� ��r�L�� ��o@f4�t��>� ����b��;��� ���/�(t)dd!�����LhK[@�e͈����w/u+˒6� ���]�����F��% 7l<h��/g�N� �Y� X�]�~�P��p:�}�5� �0d<N�;&y�k��8�(Dh�p�}�<�.r3f:)s�6� r����)�D�]`�����V8�kŎ �U���ہ:��d�H���^�
��Q@���b ~���X 8�����b�0���L�8 ����-Gn ut�����@ ���r1.���Ic�5"�S��:�?� ����	 Q�_�0ޑ�H>j�4��k^X�H% �P�V\�nx>v*��_��?��8�3@j�9 A�_[C�7�\?f��0����,��i$5,�Y3Z�A�CA�4`�D `F�W-w;eL�( �G}��d0Mp����>uJ�A Z��.��]�6����ݠ�� ��CI����t,�6	'���{�
��<FB����a\�h� ��?{|g�Y�{�Ǚ��s�0�tv �����@�&���9�J������L�ht
a���Q���-h�_cI���@?5Mvm;=s~\{ 0���Z]�B��p>H�=�&��>�~�*���) W���
- j����������B����<�5?����1���6NzsX&=��H�XJ,L4 ��� �� ��d�I8��" ^�+k��,���N�0v��>b������`�pL�C_;E�qs���2tF �+��?i7 {�.�-5 b�`����� ��1~[�A� �n?�`Y�� �Sl��
" �X��E`���'N�bF໷�	��@ ڲ����۷��H aL�oKqpJbM�vNx�I[s�$W�H�uo����%�G�T���Hw?�\�-,����Z@�/3LY �����2}8)o�\n{Uy?m 'q��ċ��,ȭ�ֳ���4���� �H����u �#x@��\ �PF�0]� ��:�Vh7% ܨ��	�� /iײ��1�RnX�D��0
�a���K�b��@م� ]���G�����s��� t�������$�f�m9Iwj��.����T��CxB7��ϰ��(���'Aj������y�c{�vB�R��� �0��`�n:6PNtmBpd�?k!�9!A|��';c~*F��s�����hTp �[���`�"� X��`�Yc 5��\�#���
�N�Z�(�0`���J�D,�|���p8hх�+�^@�jX�� �&(��g�8���x��������<_� W��ӻ!D ��v[\�So,V�=% �U�4 W�_y!���	jSMY�~��<�����������y�v� ���ClN�b'���6@���	'�ˀx7�N�O��l��#5U�qJ Z��H�K�H��D�<Z�"ՠ��	��h�|� S�"خz [u)V7Z��}�	��2e_G�w���� k�q<R�:Eu>�QmX�N�/�B�  )�����$���7`P0�h����?I�J����P ���Ć����}Qr6s8&Mx� �)�I/� ���������0��j`�h��i�$	B�y�B�W�}ű ���fuǝ���p�v37w�"yFphMst ���k��!��������A��no�|����&� ��΃� +�(Djwr�����/����� ��B2\�:� O�1u=�ώ ��J������~�����F�u���AnIe�K)x�Ļ	���������o���� ������� s��Ω̒��B �P���h �&�4�����=i)w����z$ �(��ꃡt��!;`�V�������Ӌ��}d�0�Ş�C�P�.�N�\8^ ulm������-�� �T�Ӥ�b��X;y9g�2�^#&۬= mR��I�;@�2p Y����Sm Z����PlfQ!
O���1	U��;x�P�^@B�- I�uT	:�H���h߲�utt���{���
���Tݹ��E���bZZY��J�d�鉕������F¸��ǒ���N# ��Zm0`�u��GאP=?U w$x`���^�/`)�� }v{�C9�� 	N
$3��g1PA��"� �T��= s+�w�@�c����l� k�4�I�� D�|���Zf��O���j�>`��7�W��WXa+�f������!�^��+��a�K ���:�m0�#��%q���3E�פ�z#��.�_] q�O:�x=�&��׸�aW��S@�ؕ� &�k�7���@Fx��V��@P�Q�� �E�^�� [��ޏ 
��i;v���� M��j��dI���>��8��a� ��� �l]����&�~��/~% �-�D�*�f������ gm�la���-���B9��|+�{�\���� :=�8����������X�>��9�:!+���A��mF{8�x0���p�� ��\ܼ @�v-e��D���@��*0��.L@��� ����f�y!���] �D��2�8��ɽw(ȧ��`������ Ɍ�l� �I:��O�� 1�
�t�.��@�N7�9D���(�. ��,��C& �J(�
K6
�O�8Py3�;�5�F$<=1���I ��.5�$��J2�B'�04,
��.�h�)��U9 ����
G�gȅ>�}�P A��y�1D�0>��0�T�-� X58�X�
dFz, �WԸˬ��g�x��0B&8�YN�A�y��G\��@�	�t�0W�Y٭�x�P�X�~C�!ߐ�� ,��d�xvIb��_ĭ��m!L�>C"�	L�����?����E�<�o$z���b|ɀ�;��&
�������i'ހXDB�S�d�"�"a�:T��ƒA28�WQ�۾ed��Q��+S5�(��T3Y.�H���C�����w��P�l8LL|��B	��Į�+� �FZ��D����.-�d&I���L@<T���$��d�\���M�0ϣ��"B,!��)�N���B�h�!�?��, >�?�t)(�a+����F`�	���.*P�(C�"��\�4љ��^լj��K��������,c� n��M�bt\��WP�H�|������k��߁�yy>�ؔ >IX�'L��,���5�v���=*0X�,+~7�ox��Ȉ��(܄��G��� 	�0�w��1pD��G��#<���{<��8<���Y�*؎<>/�#��(���H�>e� ����
�b�cȀjw�m׎ ��
���;� ���ѩ>��L�L4	~�	@�u �X�rQ �޵�e�T������� 
<����v14`��ʀ�JC�bn Wl��T�|��<�{�Є`�V�\���� )N_|.b� ���!��F��+��9���`���@���(nBi�v'�`D�� ��Z���B� ��*�;� M��$v��
�-`oIN+�`Z�2إ a�݀y�\"� |A�ہiDw�sڙ 7�1�h ֈ5n��J�# {��W8? ,�G�x!� ����iB�ʚc�JZ�� �h�zHe j)��+��: ��#Ù�� �[b%�}h����/*n�I�����@�Z	���owx�(�;�. h���m`!�! �{P�F�pI����c���] ��M���� �w�������˩e4[]��ThqM謰x�S�˛�k;�̧��G�P^98#t�;�H 3>�f\jِ4 ��K�V�M ��z��P� ��4������&��� ƈ(���L�����P!���xM܂Ή��FX(b�)ˀ�M� #���!�ִ%���+�ٲ*�������)�������*���Ņ${(�0J}0p� �)���2�{@� [A�uz-��4H� �ݯl��� �B���y�N�kq������%��Oz���>�a��ܡ����H�&O�2/^���#�|��uzt����NB{-^�0��k��\��8x�/�p� h�s}��@?�e���C�[�:�@p�� ��*&�F�
�?��]b.:<��V�*�B�R��z���he�'���6 ���I�do��TH2{H�N(�d�0�	��4|�6��E|��U�����~*˝�M���Tfx����T��o���?,��f�9ݏL`\��-���X�
㛖�hJ͙��J�tb7�����7��y���4�5{�9f�	�L�[01WYs4J1m6�5I�jp���n�����D����P7g$�҄)�|	{ؑ�"�D�����$�H�983��"	�D������q�K֮�D#�')���e�.����}��cs�;�5��~�m�����p*c�{���×���_�@@�a@���"���{ �)H����%&f�S���T�_
��8U�1ኝ@`���j�_(8_�u�:Rҕ�m��Fq!�8� �6V_:���~��>�� ����ٰ��[�}��v��s?ُ)(������8�y�A�\0� ��#���O�|�f��� ҏ�{x� +��*ц�� y,zǅ̍�+��X���3�#�!���O� �������� Ӆ�ɉ�Mș�(t�4Y�������z+�1��Y�)S�B� ���!��}*ˀ�O�T&���K_��x�:k�T�Y��u�t���i,s��� :8$��p�l����z� �*������jq�q��T�~#������`(��{}9璠&+��{vЏhB�s1�_6�ď�Y��H�]`<M|T@����0ރ��YM�0c�y7�1�9Y@F`s�6a���餿(��F8!ݝ�#�B�00�Q�'I��i����Tu�w����G����Z�a�1U*�{OL:X@�/�3pH~0�U	a%1=���L�XD����?�qF!(Hx���%-B5��Mt����&���\�iFp�Q|��[�"5?!�E�
x)(|!	�B|�$Aja���P�j9���(�k!TD�!ɯ��b�DPL�l��I���� ��3`!]�M��a@�k"q����ƍ@XG�@A�x�8��ݸ�H$���)��L��u�>;�֘m&=�B�<�,撉Abw$dB�D��8դ��I���$8�j�(pi��?���e ������&�9��Л�! <z���4.�8��!v��`܌ �?ኇ�����ЂF��1�.@��P{5Ȟ�I@��.\�m}:�,�a�0|z
��!�@8�X��|�&Ȁ�+ޙ`{) �� �!�X�_Ę
�%�|ā�����e�s`,�ˊ��ĉ�i}
��f�8���\���+˚�,��8@����\���Z���+*�t�s}����?֯�J`� �����!���[��� ��\�(d��$�� �3�ʪ$�L�@	��a�A*���2 Pl�|�6͎P�t����<,��k	f��&]�xTʐd�ܓ@�]X�����>�zЋ�l�Y�	�܅1���ӛv�{��� �!m9�.$���pM���c�$�~�X�41�`� ��	���z]���+t�o���͆�0��Ҏ������ ��#�{f}�$}v��:ʏ�.�`�.��O#`�įިIҺ��<�{JX�d�}!��W��@k֏���,�%t!;��lXM�� ���u�|����@��M��zW�1�P�`�����G��1�X��i�+�z��� ���,�<g�����`4u���ݵ+��\�l�������P%3����G���K�)�O|��X����!ɀ�P�J᩶1���3Ȭ�d�y!ԏ[4�@P�p���D�n ,�ߟ $��M�	��+��<��`z��4�XF�)᠁N���M����t��>��A`P�K�@�t h���̞P����} � ↤o؛2�M(��4f���(�P4�+ˉ����PȐ�, =�5��� *ˊ�.҃y� ��4�t�ͅ���-����F��!8��/���M���菶O��* `��)�����, �(���^�G������u�
z���NI���!Ά���������@�zH�\g@X�mᅴ���K�@���܌��4R��+�|��f(z�Ӆ*���XHį5�`�0*�������},AD�M�)d���4A �@��Q ͊�1���L���ɏw|��/���0}��� �H瓗LF�fD�!�@�cf�H`� )�v�u�o��7_� ����p���9+�:ē'Gz�L�`l�����Ě)�奆85̃`΀��h���L�������}��K�L8 �F�����@�] ��bM��g���KQz�л��b@�aM�H�
h�s\y��p[8u�*�HM��>D���5a|��u���&y��UV�񯵲��o�!��U��� ,�b���`��cMW�(/?"{<6`�ڹ����0f�D��>� �v��,w�07!�� ��Nl�Y.i���:�E�"�0bp�kv�0$�/,TC�F�#���Ȧ#䒎p ��Q@����i�����,�$��$�l�GQ!� R�ً�{��R��#��������zֹ�| �MB�I6�$�2����1� �
>?�s�O�"ɉ����$��A���B�BԔ��j�K���W�������E���@��+>n�]��⠐
�5h ��]Za�SR�G`j��M�΁��TU�# 1���	;b$/��;��������cJ!o�TH�|M�0��UG�C�"� g�U�����0M�Yi���4#��>QR�!ְ��c�d&�ҷD�_���>��0\�X�����[�������^нU��	��Maט�|�Yל�R瑗\���J��s	0y�`א��?T���aXd
��֕���$����UY�X�D���U���*��h��� &�ʐ^+]��g�@>�q�S栴���Q *��<7d
��\p���y4��N`���#c�� ���K��G k-����s?��\��7G�h���y�v2�o���	��k��x��74�0wF`e��`Џ�/�M�8�~bJ�l0�=�i�אx!=��	�!|�QՏ������1��2���l۱�h�� ���Z�T>\7��F�UR��n@t�U�� -%��т�q�a����( �aܹp�� �P����'awg\��\��0�>Q��y�H z-��[P�I�|?��A,�\F��:�1�g�@Ж��`�)��r�v.,0P� ��<�$��l,  5>���.s(�vF����4*�X��~�w6pGh
���U!TE�Ф� 3�Q+#V,� ���'����`	��K�tQ��9W�n}�*��h`� eJ)g�8���� �]�U98u��3�kdP���L�,�7�%@$ ��*��<y�y��'�,���>�`Ѩ�K�h J��eDE�$��dl��^F�u�Z1�c��n���@/;mI$����0�a�}��I"���>t#肐2M���He ���pE�Zd�i�@��nP�a(���Ę�,�(�� �B� ��0�:���U$�x`LX4~�*��qS�\b�	�Tp �9AWi� �m�] (�ɪ;&���?&��(l�P���qX�/P#����=<8S��X�u�bӉ��@@$��u�X=bQ������0�UE���dIAu�U �_��n 	M�c�q��<���C�s(;��)�Q��>���C��I��K1�>�0cb}n1
*�[~��0�Ǫ�e���( �GAfD5I��� Ί_�����G�YHp}o+I�P	�`蜆���$�X	cL���Yfi{_�}RG�$ȗ�&��i�����F�`x���mj
KL�����7�,�_�@�㬀MS)����X�U8D��U~�`��prVM���@�AN���� .���9{��4 ;�@�_~фO}�|� jT�E?J1�M�c��V���:����0��E璗Tb� �I�� {.rY��9в��P�`\秗F,"� �T�7W��[�r@���5��%����	�|������GDz`
��]-	B�jdz�&�h  M� ��UH�Do� �Ud-⟊�^����e*B9�|bI�p��d)�B� �[���;�FJ	�e���;���Sm��{H�1,�8U�ʜ L�"G��K�@����?� ���N���,��\n`u�e@�V� K�'��Q���Ĵ����dAH�V畗<p�N���֣�X�kO�v,���Ǘ�F��\J7� fV�[�_^td�O@nL ��+�AK|�d�h,/���᪍q�\H�$�I��A&���.�ړY�4<k"e��c�ΐ�aZ�Th� .� ��B"�=G�?ݛ����I0����G��kM�OX�	(Ds@��S甗Db� �?� ��ס��S(��  ���s�Tk죑X ^�d�.( _F�x��;�0��}���������+�CV���9I(}�xe !�7:�I%~AR��ވ�k �r���ĕĬ�\�3�n2p.kixA��1�2�,���	�&�3�H=�֕����k,Q4w����<Bl~!������>����6���Y5H.Fr�Ed�o`��4 �/��MlJ�0H�T����eyh���� f��E����B����d�����_���'�� Gx�]�����jQ�4���3���0Ot��"{���u?������m׹�����E�-dA��T!=�00rL~��q�.�F�P�B/��')M� �������<#�&���(�>�H[k*q����p� c�@�i�t4�� �/I��8*}!�0Q�(!(�{��vZ����hR�}�&�ΰ+���}��3��`A��HN`��*�[1�I0�k}4 �U��}�>+' ����\��y-�/D��]���$l@	�pr�E��`ו��z)a�G]�h���ݷՁ|� 急0M��
\���`�]�"�
`V��)����(�a �\�k�d)�����_a�h�/�;��$��,@b�g�D�`|6���	<r��cbMTD,I�D%�5L���B���; ��-�̧{1v;��`�G d�`h-t;#I�R�`.q����O�t^�  ��}����@ARP�!���*D8=�U-�p�R C��T��tp��ެ ����<R?P�Y�g�!�� @�y�>���@G���6P��{]�9�)���*.:�ւ㣬��ra P���T��ǈ�z ah����W�.���k���|)�N <\��*�.�P��Ոw��0�ܐӌaPl���ga ;��Q�M��ѳ��`0!�')�8cd���Уv�њ�؀Y{��+Jցx%�����o���ih��E7g�Q&�=*����9.� �����]\G�0 ����g�� P�ܩ���P8خ �_Tb����P1 �0ʥ����*��=!V� �K�
��������QF��`��j}?��q_�)���&����n [�0 ��m{0���٫���}(5')
8�dzx��˥��ߌD8W ӥy��Xtz#�+��|�A�����N��]D1����c�La��n���/!��P5�.���8�)ÐQ����LO�P�/�����Ł �v�`�O ��ң�� �h逐S�W�$�����(�� #����D��v��@�����Sc�����W��謰(`Kh]�u2P��xP3���g�D�h�ځ��3�-l�ҭKĀ��`̀��q&�,�e�/o7�>�$4h;����Feg�!��6, $�� ��QZH8'Y�1�Ը0P�.���Y��2r�bh���0U')��a�@��8 ���Q;�G,�$Rd���zD��ʌ��c�4�k���! ��r5aT�ѡ�}��\&]��J��`�O #$����C�0L�x���	j~#&3�!��jέ	6D���c�À����(4���D(��
|�m��vB��^ң�����f�:�o�P�h`�$�LD@���f�x�S8 �=R1� a���ze���$L��U�<:g0[XS���iP������E� �`� !"��0�����j��$�"Өo���-�pے�Q�� ��HH��7u0��I���,F�ޮ�A���GH ͸e`�� h&P?q��M0o��v�Y)� HX.����O�@�A�Ǡ��T���}�ީ��k
�qθ� 7&LRg�D>a�ܶ}[*�֔�%-��m� x|��C,lw��4�墄Ag���c��D�+ ���$��,7��O�R����W0H�/�TӨ�`�Q��� ��13��!p ����B4�R���n$/��Fp�����7�j֥�sӠ Y�*�W��&8�0���mAIɉ� ���o$~�0�+!L<�X��"�%�rd) %�&�R8=��컛��3�e�U~PDS��k0��$#�|�`�c� B��ުD�W�2��I�{���c��1 '�ճ��F3�ȕ�L�"�!٩*bt�áR��K�	 �����$m"�ά݁� l��!?�odK�@j�����P�gk��
@��ߟ�9 w�F0d�A00t�@K�!u� �1�ٻ}���ɐ���Fԥ���GdPܥ)�`�0�l:&� �TМg��Ў܈�����|{D
����s��Ee�o�X"-���0%/������r�d11D��D�M? ��K��elx����f�y[��&7�clS�,/��0ב�5)#���!z�e����c�b� %�տ	���ۂX���ʣ�����eKK	w�1[ or��$�`�8 :W���C�{�EӖAd���]"0X�~w޹���"���@$6@��&Z���N�߀�Fy���+���!����K�CT � �~q�\�l_�D�,�� e Ƴ$r$��3��9ꅌ8js~ĕ@�j�91�V��ӆil{��	7�l�@�]
i�P�G�H>������d��x�� �4�`:Ꞥp>j&��j(�;@���0��@�,��c�I3 �=t�w��DG!�܂� ��@1�	_Tj�i�P�/$`�u��K��}����¨�F�$�� ��Kd,�좨<"���Ä�1 "A��$`�	�Y�4��4̰� ��qn^���'w��|���,ޢ�����(<1)@K<j@�s��40�ϥ��?b: kץ� �1��/�Į�`e!+��x�)ۄ�*�d�ߡ��"g<]�7x8H��Q�p�(�"����dRA�[1 �A��xQ��� �P�o���6��@Dx�;�ՍP�G�B��3�jrFv"�r�
j���䀢�E�;|�\�6*����T��1.1E� tB�m;N*���S��/،�A�(���c	f�R��<�n�)�XYW�W^	��J���k}��@��/J�!<ߕ�9w��L �ۮ��?��,�$H%�:���~٫��XpU<���ې��R�薘������5���Q��@���$\�H�P��׿���Z���VI.wP�p��T��ԯ�4���Ƭ�Wlh�y��|�u���U�]�h �k0�"|(�v��������@\��n ��Uxq�� ��(!�����U�	��xDZ�,3Љ
1h ����+�^D���r������A�( �������>�.9D��yE\����+Q�FyiT�o��(��i��d�`��jp��� ?������ ��!���_$¡��ca\:H��
�䀡�����E�scT��g��@ؔ$�ь�= ��Ygi!Z'1D�����D�y�o�	ߔ�) ���	jqn�t�j���kp$����U3/�p�1	Ʃ�g�BP��b�	��e��$a=}� �7�J,m��i�!O����Ag�� 
��o&�ޫ�Q�d 4���-j"����~	aPdQ�`�fa& �b�����՘�:^?ŊvʐƳ�9�⬰@q�DOx�D��H���Y?�C���0��� o��^pN�m�|�)��#��XI艌XP�a9$�\p`߹�D�S���I�X|0&,ͥ˯/e�iե����{�
�h{�	E�VҔ\�8ۙ�߀��h�� ^~P`�,m��	�Z���% ����`�g &HCd"��(@��8:���6��呤#���͐��+e�.\#� ��Y�t�	ZWT����U̦++���T-f�����螐Hv� _�J?B���I(�j}Ĕ@�jǗd����1�X/��e�P��]K\���x�W Aj1G���x�y�t.'��VN�+`l���Q(�K�K^�WH4��ґت \Փ 	qa���d��ya9,c�L#���Ȃ�TaC����kCo����ׇ�Z���V�:�`����=�� 捫��k	��`i{pM3sC��h гJ:J�`l`�d�h��j�U�� ]�"�lW٘!EU�f�}�
��`:%���C��5��˗��U-��W�_��|�@GW����yB4�(*\Fg9#���U�bP܅a��h�q���_�q|u��`�Q3�)ehtlH4S�[Ñ�\�CS �]���%V��1�Yǅ�#��f�։��.A����� ��R�-,�J8��P�U`SX��k �Gaj�����@6R���ǆ�9|B�d%`�ո���2�a�&f���M>YU�
U����]	\s��	F�qcr�&0R��&@RkLT	��P �g�Bm�	��ŀ2J�aX+.2lP0X��HD��@P`nF���$��O�F �O�yǬن� ȀM �~��xS.���\����>?��J#���2�R�63�E:�|�C�	��C��J!���DnwV��_�����u&a��@�� 	�� -��k�Ȕ�����\���ץ� �A1؅UP1Q�9Y��L��AQ �ʆ�IG�� f��w��Mj1�"O葂sp�:*� >��P�Jë �3�	McP�K죩�GV�^kA�
�x��Q"���}�� �2��9L���@�����b =�%K "�*����R�J@��Q:���H�#�E,�o7-�@r�~��ƺ��"�����r1o1�$oub	5# tPS�8��H��)�7��`����[X�"< OF�d�RaZ�ȉT�@�BR�v�� �%H҉!����#��@��̫���۪��׃I�����P������ [�l�T����Q�S�A!��9�t\C*l N!@�[�V�j��}��;���V���,j��]2F���� ��?����y���cr��/$��n�
��m	˼�2�-)F��K�(�D�`p�5A- �Ӊ�$aZ�	0�W��)�d"��i�2��-0����X,��N%���a@RC���Z�� 11 a�M�EP�MPV��vy=�#�� z����:�s� �Y�DFC7�''V �)-�O�s:=�=χ��o���H9A��-H��$�Zm���0�И�����Ź��Y�(�ӄ�^h@<�[��L��xu�M��}��~��2��3�k��0����	��@'����;��!Q4�% �@	�i����J�U�� d�Zz�������Y�E9 �D,�� q�9�h���:v#��A��` ����i
a�*���O
��~���H��A$i~Q�&)�g	�O�&R>o$�`cA�@86݃����Z,�JBC�mPa�D"S�A8`�� o���zga�~Z<�b/��1@�V�^Ñ�t�FV ��I�_P�R�_��#64%�}mP��zA�M��P���b�f�	���\�N��%UVhR���^���.�8�Gj�v�d��E�-Gh���y���@Oha&{/���9��}Sj(V
��uu`Ah�d+��*L�օ�Lh�璀� ���~|[��U�T°��2;
C�	�qj�CG.)��(�g Eh�����}��gX(uS2`m��N��&x4�+d`��af��mQ|���trI�B)d�5	D� \�+1>F�d�%�mqAYg�	Z�!��s�"@f�P1"e'�=/+6�!`׊Z�&��� Za���D����4����%>`\�'3ېAj� BO�H�׶
93��� @?d(�?�����L���C� ,��f��9�0_��� �4��`ڟ�������G-���_�t���n�eǁ�3��Ӹ(�Ë\0U�����HO���[�s�M]Of���q|�Po��E����&���՛u�� �if�����8��� -U�q�?;X"�0�Z���䞉R�TFڵ�Ĉ�Z�� ��680J)� e&H���� �UHd ���eԅ��@�^F��_w��hXMVuPe U	EN�J/�# �̃�HR$��t�ʁ�	c��DG%�=�B�� �h�������� 6	��P-�U:���1.85�E xception9 I�f
rma(�<le�s�, �d�th��6ql�w~i~gzcdos(�~�a@d�R?�.*m� Th�k�you�
�L(fpFsbCTRL+_��6�i�md����py�li/b�ard)D6BVe�s'��=�%�C��ck*INGdOUT�Pro��[F;@�iht=r�P��GP�.-n�$�	��P"��eh%�Ð�a'$etBo��(�$���eB�U�%Cs��j!�\k!��zk!��ck!w�kk!{�r*FQ��&�}H:ʕ�e'B��Z!K��+��/��R4�(@��;���.ݡ�U���L�*4ebPs!T�X�<\�EwJ�}V��h�ͤZ�{dw2�s�EoB
iLR�)(�	���$j@�$���3xK1ȋ�(⇑����}^`2����f����=��僯jhǀ�$��% M�n!Ly�e�[�Ɠl.)���8�Y��&  ��41f��>Z�N��@S{8.�P�KK�D��t|�:zp�0
a	\�R{f㟬���i�$�"�`�& _��@w�~���ev5���`X�h����r����9�e ���A�������P�._	@ɹX7�>!��5��`�x��n��,�� �I��Aw�8`�)Sp9>�R �u���Q�!��a��V_d��7�@��>�R9�Hސ(X<GC�Q�P����I�!���gXZ~�Q0<c[98A~BP��a�9�:��b�T�tM`�#ΰ��\ �j���/� u֠�]��+Oz�! E���w#g79P>���O� �WZ��Q��� ��<���Ф^ƅHO� U��|��>��y�L&��_��R�#��H�W���bP��y� Vd�kZP�0�5HR{4�v  �u��t�_ٔ�c�!k�[q�I�VZ�����EPe=0:q�|����%���ra��09S��8 U#(="��d$@�@�\�T6�^d.@�#�u' �f[s<�T���߻�����F�� M��'@�gg�y�O�0<2?F���8$���,D�u(����	/j���� ��z7�p��mH䰉�"z�(��"�_�l�c����$���Q`��� !��V���0���9���@d0q u�h��C��w�v]bl�ZA0�	��d|�09�i������n� (�):W� ��XF��')���h(\p���
�ǭ+,�
�f���k!��Y�ad��crT?Xƈ���J�"���Re��a@�1��NY�T;͊0feХO� �v.�}���w�Y�@*����U������8�ܘ�l(x+4�S��X�:���J �9:��w�,?�c0�n U�A��y�X�xu�p�<��������É�Q���1#�����M��>�0�O�AL�x;�v0��T�,�3�R��0��0�����j���>�1fOH���� ��uσ$�)�>�@�bܝ��y田"���[� H�9&u�\���{=�J�p.�n G�B��BLd�$�<��n�d;�F��׳$�:0�����fU-��I� 9���R�2�})�@㉬�[�;�0�W�>� '�O���c ���ż�b ���ƽ�I ֜�U
@o����$Hg��(i�>B �J��x��yu #��	�@� =щ�gV���0#��`	��i@XȈ��+�E�K� RF�� ���dMQ� ��v2eB�����z��� ʑ��!~w�	��]
 ���U Ն�����j �mŷ0�H_`�A��3��L ��F �J� �ma2WH7�eM��<0�s�� �r��2����W�^
�q� |��ӷx, �n�u���k ����9�28��У �o�6r�S� (��wp��䍽�P�0�W�NK�(B\����#x� A��Y��F[���U&v�:�d G�P��(_�2O�� >�:a� ��g���� ������~ �ڕ�H�m� �-��E�k� �#�ju|�P��@�;��$E�y����` 	�Y׈�����;�D��x�-����� ,<B:�X�Ajڪ�(�����._@�7m�a; Z�R29]��ID�9 1�X�uJ�(X�W G�V���� I�O����% ��r71��w� ��)FiH�@ ����<\PW��p2 ��&X�F��� ���R����o��P ���b4��;��@a�"�$$� ӵ�(R ܞ���*K ץ�����$	?D3`�Bz *%�6<�LcW�@4��۔ x��N����	�(;i ����m<�L,��H�ך8h(�V�� �����bo�hx@�`�@�� AI,xb�"�)m�`J��¢�M� k\���y�� (��Lo}Hu� z鰄�%?��} ���h�Պ N�@�B�Z�0m8/1��_�T�NR����+0��;X<@Ԩ8���t w�,��:� {�*��9� v�(��l� �G��j� �F�~g���I�!���R����גS�0`[� �/��o��t� ����s�� ��,$�%� #΅"j@3`�Lc O��t�� �fy�R8<��g����� q��x�ڡ ���!�� ����\� Hp�gQ���9�!N�F3 �XhA74r�v!o=`�X@\�Bn
�����XL= ��?��� � ���d��Y���or����\E l�eR� �����{�w��	'Ҧ�E.]�g ���*IZl8�V �ɋ�v��� �-[��q}t� 6lz�~� ��Y��|2u� 3;���c>�4�[ R�p*� �,7{�'����^A��p ��`��Į ]S����?<�X��I}_OV�( ����R��p �]�Z�0 j�J�y�^� ��[�?9ʝ�����,kj�uȀ���G#wA�@�`� ;��F�Uzg 1S��I:H��a�{p�N~4 S�#KR��G}W���v)���0� K�y[6���|	���] P��D���	솵����> 7(�S���9w a: ��JV���0�İ Z���	s�� ���e_
 �9I>1��� �U�3#�O�C����($<�� ��� ;�맵j�������)UTL�`ݚ��R��0}��H/�� �;� 0o72� !3l<;
��n� Y�ں� �hė׵� �\{���,�9�v���Q򟕪�|�]
��z �NLG��* �_Ĉ%W ����d �VX�a�Z�*��>�d"x��e'���s�w@���t� �����}s��*���q�����:�Β[���,HxP ��X� �G�ؗ�(�H� ט�)��O�!���֝�1S�ܯXa���cw3e��x� U�����h�����\v���"��7�P�Б� �;^������aT�@���uo	�}DW ,���w �X��v�8�x�0�w9�:�}G�дv����wX 9��M`'�u ASZ��(����%�8<`f P['ו���gz]9-Q���V �x+��(d�)!��d����U� gȲ���c�mʫ�ŀ]�k7�)$�`U+& "'�E�*#VS>O�<@3�H�����{,@O�L������������C
6%�0lY ��߉�Ճq����#p ��v�����@V}� ��%L��!�e�);�+U�9���� ��;l	Z��(��c�L<�ӂ�ȈO I=q��)2���j� jr��p 9�۽IT �-O�=6�" 3f�ϙ�� _+�#�-� ��G\�Hb���e#�;�Kj2AM�4�� �S�]s�<$�X< ��߯Q����. �O��ާ� �*�
8�)�P�Ί .�[��& _H �O�p��J� �%9VI�P��
wX:/. Z������ �zO֎w���( I�Ö�N���S�2�~��{F�=���d��+��|�023Y]�8���)��r�u(�{��9� Tk��wq5 @2e��ڦ�\�3.+���) -�ˣ���&�(�8�����	i�#S69�� �ȍ�Ӧ����N@��]�qs���>��d'�����"�a��fzϖ�v�-!�=yH /�,Q��_� �^;$`�C��XÄp�$7�H짙d��j�O�4��2 (��L �eM��t`�Qʨ�� S^�G��� 9s
Z.5�L�4'"�7�`�¿�e�`.Z ����� ��v"1g �u�,[��fh/@�������G �X�/[_Z
��J�>����c` ���V��u@���\���T��Z�Eہl�b;��N a�_<8����x~}���Ԫ1H]	Ȥ�`*�#N��<'���KzA�Ӎ�J��|.^� ��V_���E Վ�S���:��H, "�H�*O B�����A�9��?/����E�L>Kx~ ����=�)k0t�`����x��0����k�@�(@�UnAO ����h�+xd@?��{� ��|o������u~�@P�C��O*���8�����s<��b ˀD��_^��p8� bS��L9Z ����j
� �x��g��L�Wn��D �\����/^]"��˪���.� ����[��� #���`	(�����|���$`� �����3�Y��ˍ���+��6$,�� ���=9��Y�}��;j���5�� �c��?,#�� ������% ���VAU.�0 ;`�-��P���(C}�J�:��$v� �h~A�>�Rm�a �,Z� Ѓ1��bg��~>��(f�5� ���&�����+��*��tPl�
��[�4�8k +u���W�Уo��N����r}�!�h��CmE	k��d�4�Ćq������L5 �K�!GW�ؼ���,� A���U� |u�}���VJ�#6 P�;��q5� �T��>n�Vߝ{?���`+v �~Sgt"c%(oh��w�Q�dE`�U�c�88�����#����`�n�W� �Ԁ���� R��]�*<M ��y$=K�� ���`�
d���h9�0w�7	����Z��R$xS�%M�sJ�O�Ѱ��?�� |��)k-��
��@�� �3��Ǳ<��8�z��X�p� �:���B3`x���j`�<�> t�1h�z ��b��o��w"�U ���n�^��Y`��#b& O�e�I��f��`AL�{�����+�ȠU\ �G^��k ��m�l�Y�]$���� n�H�SV�� 9�&%��� 7�,+�#�Kl�f�Z�b�j����]�k���h�� N���[J�{� ZKM'6b�) ��V҇�T� #�.�<YAC�H�ܠ\�	��k� l�E%6,S��� p�U��jP���mAH@A�c�*%��Tg9<��f�DT�,~ �H|j�@�QXK\P��,�W` �z�8'χ���d3���k����xw�@����x�cW���4!Y���N�1����߄&� ~*�U� �[L�kP�?N�"�;w���v��c[ �����(�G�g ~�䫅�� ���}�e�� *~�I@ �z����w9L��U��cHJ�;�d�� ���GgO�� ��X��+wjШ��?WPuE�# f�C,���c:u'"8�	��VD�a���e�a,�����( ~T���"O���=&��8)�c1I�0�h�W6 �*F�2�� :OSz8X�������f�g�����&��߀Z�n yO<��7��	�^u� ���0�� C\ ��`j}:bf�R��. rA#�|�p2��9��-�&�I�n�f�X�Hմ�91 g�q��B<�@ V�{�_fm���>5�)����̮cu �p(�IW v����ؾ 8��g�r�. 6��~(�X$�n�5���x0J[��w14p�K�%u,���ā 5��ǫ�Y����{�d')�!�o��*��Dt�D��D,��"�s")�"�aBlCe!L�Bx)~!Ob"T"�|B}�T!`�y�Y�U�<�ODE!mH������J�$+C��@�6D�A��+ >Ӛ�� Z��?�E�YȨ�C� 6��ΰm��$�s@��@ �<��Q�L^�����F�%�1v���0@ŠI� _���:�E�~h��12�����}a�@¸)ģ�~1pj)� �L��}$��pFN��9��E ���:�;���!�IR�T�'�1� �^;Or�P���э7�)��Lň�;�hǖ�`]<���(����Y-4�X��� ̚ ^Ō�5� }���H� >�8�0�1��$G����7 U=A΀]V+�l� R�c�i���� S(�d�j�zU	  ��~^��/G w�Y3�b� m���~�h,��� ���A�
:�U� p�Z�@�>� ��Ŕ�3� P�˳���}l�Z�L�dƐ.�iv[�_T�T�� ��b/�:=�� (P��* �Ӿ|ޱ}s :k�����X�I����0��u=�L3c��5���f�M�4�P�����# �s�&�o�?~Z�� T�A�����|֎�9�瀬�4݌���s�1㎮��v�4ɐ��!�Wހ^�k�Z� G�D�j�� ����]��< ��7�o��2�0ـ�U$Ъ,�տ���R�%. [�z�@;j�`���I>�Kē�5�%  e
�s�� w�F"�1?,��J��hD�����P��6�&� `�����W�s��,���.��T�� �8�| �9��0݁\������o��.�4@ h���LJ�:��C���=�e �|К�hҖ����G���B̀�29gsg{��0�t��R_�>r�@��:�5#����= hj�۔䷢�� ������	��H�oz�c� 3�pE�)����S�����݃�{ L���}x8E�� [C��byA �	��i6� ��]A� m�/�e�c� E�S�s3� �.R)�n�u+<L
0&){p���W����4�5y ���Ғ�O ~	��!���m+z ��:��=��& �h� �`�:섮�/	�޴� �b߷f6I�AбR �� ubw�4 CŢ(%à0^�u[s��8�ҏ: �G��#2:�Y��&��<*, �١��v� ��Q�X���˒�'p�S�r> ���N�`�:5����r^�ȺZ	 W�/���@� �()�EjG� �����L� �J��-#U�Lj) �p.��R ;w�`�(2 �ULf��� ����9�^��@�?��ͫ.>�,�@n�G�8�m�^�H��r �Y�Q� �2�yi��n����FE�k@ת�>&�DN ��!��\��b�y�>� ��mD�V��t� �n���_�` �s�:m� A
k�b#� \}���� :�H��� &�[�!��� h *�.p� v)
�2��DSF  ��� �z�<Nv �U�%�F��r�|����0D�3��������)w��[Zī`I�8 �D"���u ���i�I�q�v  W,�9���V�� �Z��� #<�R�� ,9�V�JJs@�?��,À��5o�$-� �e�j����v�`�i Gq��o 6�k� �`3�/�n i�m�� V=����e���cՏ� n�Y:l��% �m�S�M�� �u*�|�%rBo�q$"@�A� 7�C8�� ]�|�P�	�Te�$�g�?8� �M� ���x�.6	DX�Y4��� �[5S�N ����tp� <�q���l�cjV`=��x� 3n�
�H�&,�� P%�����$�"�ab�9c�Lt)��O���N�� e1Kx#6u$o^4 ��"�S� �L�}�M�� e�.:�a� T������ ��G$�;��T�F����1 �Z�����.F��D&��0J;P��Q օ���_�y��.�R�@�� %�P�F���+�Vƭp�GY}��Lb��>.@�Ɉa��鮙���g	�q"�N��?=Y�� `�Ǚz�-�?�b�@ �+0%2�vw d��ne�l#c���Xu{�9 ��P�H�U j����> �T�J�� C�	A�k (7��H�6o Efm��O���J_��� �%�ǗM~�p�c ���[ҷ�!�{���`bC��L�T��&�>��`:�Kg5� Jo�P-����A �M ���Иx=_��#��u�`�LG� p�_�I/�	 Ҩ�Z�A�?X�� S�D�@��,]�|����6�@��|�!"zġ�� �׫+ҥ�	H��Z�$�艞x� ux��:�Or����j#�Yi��� I3�B�[Ϳ�w���<��|�J���T� ���ɚ������;����d���v+q� -N[7�xȕ ܾߺ&� �`����j�mx��X́� ��_�Y���	<��a�� 9���K�̮6�T�	�*���	�'Bϖ��r�y �A�]̬@r� ���+�m� ���Y2g3�j	�z�D� �TMd�-'��(A�h��2 ^r65�H�YI�����\�N�b�E� jՇ�� ��`�j�g�$�� �� �>4�L�2�0�`��??�>] C�J�LH� t#u��x ɿ�W�NѺ ��V����1 *E('��� =3���l��=���� 0n�%i���f�8ʸ�� I�����
 7y��� �B�����L��y.��� �O�A� �*�\�B� ���4�9Z x�5�m�� ��ʈ* �@y�|��� R/vh�=�j�N@׈՘��욪f�@� H�P�����^���7���g�a@K} ���Q���2"�R���� ����n�E������^��A�t�
��X�`<Ӷ ����P_= <����>�H�X�L�î D��`T�|�ph��s�_ ~���!��	йH� w��h9b5��O�SȀ��p!��@�x���`��<��"ϊz��b���gY�����q���0�< ��C6Z��:
s�mb~��D���t�Z� [�l�G���H�B4��U�n�1 ӄD�k�:� X����� S��1Q� �;ׂ�EU� � B��@� ����*H.�s����L�C����	U���j"-�`7��k�,;|4 `ـ�
� #�=��vL� �*�`Ҡ�q p"C�FΩ�(SO�/�u� l���}>� ��Q �G;) \I!u����Xi��x�U����y>@@�+9w���=�N! �a��_� ���Wim� fСھ�Y�F��L�F {p�x>� 5�d�	'u����b� ���}D�z ��gM<ʋt�{��P���79�� �d�=�fM-��,�)�E ��[ ��^�୒�"�c�Fݲ���w��Q �K�]�R�?y[� ���e��� 	����@X� =5x�Gy�I� �q�'�i �u^R�v�QU��� ��*� ���Y��� <�F�cgO� �~�M���l�/����`7M�����h�k �Qe��6� �����,G�	w�2"��/\�� �Oe@�'*�� �� �f)s ���%~�E!|��2�(�:-~�)p�I�T�t�7��U�b�⏂�S@C؟^) �e�L��5p���8�`�8X���Rn@�{ CeM!�0a>|���y)�lܵ!g?ʨ��ݮ� F"S��Zs� }瀴��E� ��nַ�l (|�	~T!2e.�k���+�Q�3���$������Ԩ\| ꤕ"l�n�d-���X �]p�m��skڪ� q�O��� ��8��θ� 3�C!0��W��/+�(�+ V#�~$2%��,@ � Ю`�:��N�՗�\, x��cp>1дꭃ��T�6�N�` ���g��v� &��%� m9�n���z͟�Lx�{J Q���ʛ�,DU�� ��@ǘ��x EL�&5�;��� !����g,%2�= #5��6G�)+�����J� �O0�~��:^�v_�CϠ�G�&���ۀ��1:�	 d����9~ ��2�u+�=�-�s�.� '���by� @�?�6��Z� �هC�7ۆ@��{� �h�-��w ⇢"�/���j帶������,���%0� ����n�7��$�����.h=t�>�m�ӗHd�Xl �V�C�) ��0�j.�	w>>"���T�~q�,u�5�dp�� (�d�p�)��&.G�qe ��|cJa� ���±T�{ y��ȡ�8H�B�����n5��#��lC~�
␀��#� ,*���c)�K@t�2�:�Yrգ  �o`�Py�<T�\��Ɵ�¥�  �r*�)��ˡ��qc �t��Gk� �+"�D�L Pd<��ڻ 1�v���O  Z?gal�Yu� ���ne�����I;� �ة�i�- q��M@w*?7�z�� p8��� r�D�_y�R K�c֐�z���W�8� p��z_ �D�1�H�ΐ\ �����N�2�QH�7 �m���B�`�U���J��`�1V��l�Z��OU�_C����
 ����̼��~ �V�֤�3Y �P"�_��u.+�}�t��t�[ϕ��Ԑ:ÿ��Ҿ����{O,�k�S��=�.x.� �!�|ÒF�]>����Y� �����^N �6ˎ�$�<�iL{ `�|�4��|�vi���ܑ�� �#�w���[ �p�2ޏʇ @����Cr� �T=[�F��9�̀4ԏ2���la��N5� ��d	q�e� �+Ь"$��X��lh���(O4� ���Sh���������Z��N��Y{#k@�\��l�@H� �O^z����l� �H��#�\� !���_LP� <.�oy��?�F�J2�X�8�\���L�D�*U�xu ��޶iT�˫�=(!P~��.��v �0��q��p� !d�:�&8��pmS3��}�?�B��ܰ �G�V�u��i�cN |0m���n2�]��K�����z �V���b��>ĳX�?y ɖ- �3�~�|^�d�N@ђ�'7�Tpq��z:�da����xk�T� �0�e�ds���Q�U�:M�o$_~�O�'~��	��� etk��z�!8�'$�\H��/G����Jׅ��б� �P(t�?� =�j��^ɡ�����~��59�F� 8�M�#1���Y���8�Ed Q�J������ ��M'�bv��i� ]�,S*}U��t���N�Iùe�\�W�h���� Vu��i $N暳L����?�X���m�i��(� �M�Y=5H`O��@�30�@)C�{�a(�=��క�� �9�,�D �[��n��>�Z>F�?D� �����1��U���f������M�;�tl g~�0r�N����eZ�� |��JnYs�j��@,e�MX��nj���^�=�\�<�L*hD����1�`�v�0�
ࠚ� �T����p̫	!`�.�� �ta
H&x�L�? ���K�1ʷ��q| ғ��ǒ� ]�u�S#�� V2&�_�G� �|���.�AZz�!�в� �`�o�)�r��\�@�['�qC��K^<z�Z��L��w�
͌�m�b4x���u kI���;F��Q�=���0�	�{()�4��;<��JQ`�鼠�9�d�F0�W޸ �>Ƹ�d���~F㈽�]>Xy �2A��q�I��ɯ�|-v'�@�� ۠zE�[��0�L�@ �p�ٕ|����}�	r�\�*�C�,9�c�f�'� Ht���e! �B����	�8-˽Y��:����/� �J����*��^�����ǉ���H�� o�"ƅ�I� D�����x� UC�Sz�
;Ҟ غ�`&y �Yc��.�,ӑ@6���W�<��&&� ʪ��F"w�Iˀơ�R��' @��g�o`�H���a���k_?a��V-��� ��Th�� �I,�m�#�f�b�$�kj�g��1t�"��e�d Hg*�]�s�ˌV� �@x+P��R(��yd0� j�<wg�_�	�ۓ�`җ�]V�� s
BW���� З�;!z�H#�S��{ H� �Y¸B��z���D��rg�)��+ٞ�y� p)ԍ屢�6�<}$��`da�:X��>� F	ZW@�v]Y��{����(Q3�V��<9	�#B���
�� TI�9+ 1�W����	��b��[�f ���Y���̖�޾�68	�!�'����l���Kv)�	`����9�,�k=X, ��<=�4 9��h���Q�R$��̳�TYŔx�&�n��i����܀�=�M&��Ā���"�� d�/N>��0sg����t�W�L�=rIj؊�� I��,r
�4��� ��@Q+�`@�@���-Հ�QZ�x���"��`�UeN���C��~��3u���h. ��-�2�jca8Pxr���8�'A�*D�oi4�&ٺ�����D ��Z�k�vq�y�X{ ���R��:o ���|v�N���Z���V�	��	�Y�A! �qld&�����u��`�5X���(0eΙ��Y�P�~d��4��x 㞥e�*�%�L:�!��� uOax�rt��	�)C��d�6q�47ܼ4��r�TA�@�s�ղ���YJߓ���X>*�P��`��Ә�6Y��d`�Wrk�	v*  {��b7 �P��Hi�l��Dp����?8\�C/�����&m,@���C`�̹z&`o!�4��0� )��Dd�� m�C���=��:�!e�(Pk��v�f�t�	�j��@t� !���-> �9�7�0"� j��E(!�� D�Ytl����)@#��(H� �?y���x��[ƀ�U�DCe��.��� ^y����ϯ�KCy�8�ٖy���æY[���< |���������[�8���d�f(�w�� @5E��'�* d�Ѱw[���I7ó%����o;f��g�)'� ��>��vX
�����<V8}�]0��h�0�N������K���u��8t�{�/މ���D�\�T�f�B��L6J8��1��pNfC��a�$9{�X����k?"��m� y9c��>�˾�ӈ�]��Ԙ �F���!��-,(�<{�p2��� ��V�Yr� �\HQ�2�}��PuA U���Ώ�9�G H+�����ȿ�Zx��z d?��� kB�Ϲ�C� �����}� ��5v�t�e�a۱��s��1(��6r�<���G��0�81� :�5�����7ɖ'��R�־Ŕ�� x���^� �3ߊ�:�v� �r���#�c�[���
a5�0Lz ���p(�y �#�{�<x �!����;��(�<��%�y\��nʈmq�(�{ &�ևkR5 i\��D L���� �@�:�a������&R�X�`\����@$��c���g�
�OضO��L���m�5h���N?>��-q� ģ糼�b�]^�����D�1� x�ӿ'�Ԫ0ؙ�Pz%�9 ٹ�Jk�` 	!�i�2v� ��$�F���5N4���j� ��_tשR�~� @d*\ طb��R� ��n�
 �%�N���� ��L�u ݭ2��{d ܃	�x5�>��z��� �6�:n����Ap%��*Y>n�E�]�|��*��K�%>�=���2�@����[��M�p�d�5٩8 L9��$�.�H }�RNk�,�Ѐ�`5� �#����:�j� !�_l$�V�i@S+�YB��/!�d����p� ]  N'_��d��A�l��#\ -�;@�J���� x?����d� D�Ś�M���(5�,@��<�\Oq�̀ Xg��vW?��B�F°7�f� �Y��%=�ɨ��j�P �:?��= �[�pj�t��DE����F ��_��*\k,¸��?x�+ ��2@m�H�$�y�f��@�|����ڦ�_� ��I�?�O�e�� X=ּ�1�:��	uON��E��� ����d�r�Ҋ�,R�<���S*�, �|�u/U&:���pT	0��4��򀁷ǘr��l�n����G�1J��a B��/q��O��j�`,� ?�����>@�O9as5�W����d�$��P�I) ��l:��s��V����$���et� �Q_���o	k\���:�0iI^!�$Q�@$����yj�L�x Hg.u�o����C�B)�r��1�k�o��+ �a�h ��^~�ϖ �T������X�o%)��C�g�b�|�� ���$�� �ىx�,<��p�Nd�\J �8x�U�{�P��D����p�� ����?�rS ^��Ǘ� �ܽ#RX� Q'}�n�Wx �Eq�	��	���[VH��}�?���X�>^��(�4% L��B5�w�|��D" �z��� f�7���� -d6T��� W{�~���0 4�e�d o���x�H%� �4�V�C�.=��X�F�@o@Pb�Ui�k̀�N"~ �l�I_�R#�m	Fe�d���SpO=���娅��'���˥�	�`w0 �Ku�)������t��3�r 	��E��÷ �/ŋ�H�Ol���Ր���j`�Z:_�XCr����j8����o�`�� u�_.��c� zO�x�����8����,� w����%�_рx��rck�+��#��<段X�b(� ����]��P/������� ��U�y��p�'��B�G ���%	�#�����5�����Ǎ�8 ��`%2'Q��� ��/�!�H n����� 1p����,��! :�d=�@ �9��п'  NΓ�A�`x� 7�֤L�2 �DQ�d!�s�`+���H� -�ҩ)�� u���Z�� -撀U�nꆏ�� 8�N�a��zP$�����t �0��o,�:�_�$몊Y!��xn=W� ���C#�� >Mx�Z� e<�w+\wY�� E��'��ȯ|`̀<I�;�>�m�T�2�x�5 ����Am������F�4P-���H�/�0���J$�RЅ
pɜ���~m� ��n�B!��wU`V� �9�O�9�<�FX� 1:k�B�]{� ��C����h	�PԘ�r ��W7:�] J (�}ǒ���� L�=�kԙ�UK��Q��chOB���԰�A�C��`c��iǗ@�%kL��&c����ݬh�E� ;ϭ�W�@� <��I�}2D�'�/���uT�A��I�
�<}��J 4Զ�� ݹml�{hIt �<�z���J��n D"3f�4�� D�dr颊�:ۃ ~�\��� ��j%4x�:v�����A��(T�� ��Ie��0 P/j�������+Ǡ{F��҂ �}E��(�|����l�t�0�)�����xw�� \�rXZ��_��@y��%t�
%��`���<�~���=n{�j-���y�5)\ ��w�B' �^��g� غ�Rֈ�� 7pX�W
'y����@�/@5 ��\fB� ��'݄�1� ��:��� ]��;�	�z<<
� �U�F�_�.y� ~Yv͘�� �;:����� �Y9o���\ޛ��g@�ݓ� o���M��=���>���އ@��ܞ�h�E�zҘP�@�|�O�R��T	�w�z[�Tv �ـ�z���%���� >؁�i�� ѳO�I�S� ��Q�b�-t]��:�0o8 ��q��= �ŒD��,/�b �<� '�����W�L����R�\�0,G'w�6Z�n�Xc
�H��9�C���2�B�k�4(N0�/	�,r��̐������5]ċ���� ᐨ� �t �3%�2�� �!4�� N��@�Jd�1��T�h�(�Q�]j�,g ��`�.Hs� ���%�\f� ����B�� '��A���� 6�L�>�Y�^G��@� 0�J@W�q�:[��L���?�
�H��Ї����f���a��M���v�VH)� �!��� ��L���F5ƨ;��=�%��E�����9�	�R-�� ^�bЛ���_ P�QJ*�9� ��H���e�E�U`4�`��΋$	w?$; ���/!0�N���$5; H�^wW&3Xߕz� '.�2�y�`[�Ar`̼J�juR�W��?���!�H�Ӱ|�S�� ���Cջ��� �]��320���p�(Ή�>��}�� SAܣj�: 1�
���� X8���?�h !et��� l�C$q�D�&�o� �햲f�
�{W6�|�o ���p�i�x'>X@�Dq�$ˎx�7ᙟ��"�y��f}� R�|�� w���',lH��Z ,�&x �-�ڎ����	�"W$t` ��b�7	w�mJq�x`��[p�j���l�f���:��� �1A������ ���s)�� T]�:7Y*��@l���C�LB �<��8�&�y+ x�P� ��_)]�K <�Ν����*�4[���W ��M � ��Z\-.�N� 1��� �b�f:��ҼC$8�H�ԭƐ$ ���砷���@����� �.r�D�J *g�E�] +�'�[�|��M캀ƫc; y�a�A�F�>�� 3q�	�G"��� �S9[:�x�"���̆�=�����iz ϡ�� N�^�2��'�mh\  誎�	;�Hgp|�k�bl��O��]���J��8C��޷����Ѐ?�9� � ?�E4�6� ��D�Z�% �]o���" ���2�3 <��:��i�'��hh�H� 8��o`M,y������Q���	��`Ա{� ����).��
�j���<�ܸ����c� eg�4�� ��م�UD����pbP��. %���m� r��y�b�7_g��T(<ߔ� �Nz�ݞ��\���F�Pur�*�, M-'��$#�%�2 `�ۤ�0.� �٥,��#/�ĉ�r�Qv& 3f��Xwg�^d,d��u��� |���YH�2R��G�nx�2�4�l�$�\� bi&����;���(`��+ _���=��`j �B!���X�;Ԩ�蟨(���`�X����㷠|7n�Ku��xY�*�l}o�d�?|>�h�m�&Y�0'.d@�p �� GK�J`6�����%$؈�� �����<�|����D�0 �O{�SR�d^f��9al`&�����:�@&br ��Z%k�g�0�B�l
�H������ ���:�K"~L�~<0 ْ�gጇG ��O9���^�p�d
�w� z�iy�c����`�T��h+�3�9i� �4���Ll��2 ���4�k��1/���;�Jn�`�F�@������ ���c�E[^� �I������,X �īã���R3=�_.����S����{(� �V$c�֛3P��!��P�-���
�;/�@��8��xFX�7x�6��	�$�׼��� �o�;n۠��k S�h�$�q������Zx� �W�}��3�  ������� ����}���� ߽c�Ө�;Z���TrSL��Y ���ж�W��1 )!~�|\��=��A��*D���&��n ��e2��L �BQX����'@�L��E�H�n��� �$�PI�D[x�e:���@�
V+GD��Ja	��� 4x�� 4PT��l�$|�> ��E�!��.��t����ێQ�@�t.k� �x�b<������e74�ͧ��<3 b��D�®� 廂dI��! ~��Mt f/�;r��"&_5�:�^P��L ��ɘ�� ��57�(� ��U��{LWtg@h` �>�
�x�?ѱ~	 �Y�c� �����P�gII/3 ���`OVa ����n|u��d0^ ���������T[n1�*덀��d��C��A�+}� �6	aXҹ4x�hJ9y��KD�' ���/e`3 O��G�$�Fx�E(�����@u�% Ne���{i >;fcqg(�bl)҆�_�� o��KW	d�%��|����B�G4K �:�M@7�!ԡ����K�&�0�A�c$j*� I�T�0X� �l����vP�I9ӒυX��c}��%�{�����Ҏ��\t�v7�Y�F�#gR�V)[��|Y+�Ae&a%0�C��i��^w3���Jc�(E!�x��Ҭ��FH!9����v��~�%]�90��q�
C�N�D6ו��_|�j�=	`&!�f
��:�|�ӻP�m+W`(����N��`Ւ�V�aQ\e�����wV[�&z��8�E^A�@f��<��E�2����&�<U`e.��)`��a3a�Y�>@t�j�d&zH r��9����x/\܃����`�]q�L)`Y#�
��?Ԍ��A� �}.��9�(�� ڽ]f0K}�ܧӜ�a~S%H�諑(�RՀ{*�ܘȐ��j肃�SN��6��9�$��x���� yf��j
<�����O-�1ӡ�����V	��$A� þ;ٕ8v�*�[�7TQ��_<��x�Қ�Q$�Pȁ�I{�����"=���x
i�[�*@S`�d��3YH�|
}��$"# Wd��o�T�H��;z
���$�Yb�MN��R��p��`#��c5���1/��m�AL�
�<���gU���^q�@�(�x��DC�׻� >���6� $�i$D�K��ӱ� ���N�ʝ
��Ж������JL��#j�w�0bB#����./ 1�g��۴&�� *�a;�ꮩks^�N�����g!�>�ф*0��¼0�E]^��"��E�#W) (�� :�gj� �����@��SJR�@�L���-���Ĺ�ez0*%8��p`��N�|1{�?�k�`�]�되÷MA3�j���9��V$�1 , ��Mg�9=Tь�ꤙ� �f�O(�|ej^x}x�$%7�^F*/��VT^�QT��a���^�a�@�w���[�$`� �g�cWQx�� ��@Qj����i�� ���Q<HvE���"�v-#�Pz,i�p�M� <�o��Sja9>���x�t2~���9�	]�H�� ^y�ʲh$�@�@X
�`yq�x�'Q ��mA�~NF�E $����T�� �t�r7�~��a+�If�Fy�Eg^�G��afVr�(�����N��xF�Eb^�g� �E�ߟt6	�"��:��@/�� ���TZ��ɠ���Ȫh=�� G	�R� z�8r����&���
�Y�w�Lh��<���0�V�	fl�
��j>�ru�t�E�ȅ��f� Ο�����GQI����. Ep^��@�EDu*,��#��<��҉�@D)`q~��� }�fG�9H�Ђ���!��E�� RJK�4,l�lEUDzBL������k�) we�ϒ�2 ��M�O�D
��l%�ڄҲ���\�X7$�G����j��>Za(cb	��1�` �l�`F�d 	�W߄�V+^�O�\ �!sѰ����׈4��jO3C1ц�D:?�-�5�7e8B<�9�n{�<s;HEd�0>�"� �Xz1r�: �D,	��8CF/JH6��f3�=0�ʩ 2�Dv5�7-�/Qd���������d�q8< #�.{�+<���u
 �iF�Έ@��Z�xk�a�x\��A�5��f�/��zd��Q�A���B`#�����9ҏ�<�<��g޶+ ��AswQ��R���y0x?��'�ݘ�|%��&0���)0��ȣc���9����r$���0lз�hhg-Ф
Q��� �P�� �	�[��wl͸�@�~*��]���B�	�W��U��So����A w
� �:�	�dH�0VF  �?�VO������=�2~� a*<^��bxi��Z, 
����/���?��#�L Fl8�0;' �b��יH�&O0b=𗚀H�8,o��3���;�H�@�����u�A58� <͝��#���^	�ԧ1$����̲�;0�> �����m8l�@�=�3 ������
��I��`�y
�#�C?DZaq82�'��栌�W���@&kO^3(KJ!�jY�yB��.�TMe�DHy sG���_w� ��٠V�[zq=�(�F�-_��<lR1�3������|���CMEPw��@!<�\}��� 1A��w�_����ə�0���N���M��O.�#9 Ab��|���&��H�B�7�}a���9)�D�"�5���M1  � ��ƣ����Դ^J&�����\�O�L��(�X5��� ʿ��f)�;�. ��o��0y�	T^A#PV�IJ��,6H�G������*@ԋ��i� v�����?W(���VSa	���6��(ZO�lMH �\�T	Z$���\M�u0,�h���pl�@ �ڛ��hy	�a�ԅ�27�L�*���ʳq�n��Fٿ0H��U�a���\8� ���d���jV��� λ���
=E��d(\���8������) �-��C)�X� g	4	�1hJ�b���L�>��0�AČG����$M-?4D�B�tS��^�/�R�U���}
�c�D!��Ę[�~.�����גQ���غ�9���nA e���7U�1�_m��\>�B�9P1�8����������l��� hD-F�N�
���ՀOg��`�h�0 �G[�4�D�C�9���%%{@ӕ��P����lTm��%^E�e�,�O�#L�i��3[��d;�ϗr�w��ƫ?l�PR�>�H%.4e|�ĉNw �|�s��%�M�lˁ����>�H؝Ԡ��[�B �;q��0= �2�����R����c1��v�$��X���PWÂ���"l����H���9���4�d�(@��H��s��G&�k��4����yB4�T�  p�/��p�Q��/0���Hk	���j�c�L��aa�]J&�:qM�`̘l�+�Ǿ�%�	�2 �(WNN�Έ����!�d)�]��1��<��b �SC@��˕.~^d��� ��,��"0L2�(&��<�촀0�����vm���/\ �i�ެ �.�
���Rj��vV�����ߌ~ebgX�6����z?b fX�)����5WO�[Ć�( ��o.��{E�#Є��i�.|�&��Ea^�+-`̜Ev
�Y���1� �r�SY߾��'=��|f���&�/Qq*^?`_��tl(�ݑz���AP�@����@�I�ˢ��ax�����X��Y#S\�P�r��� nI�Z
ڎ	x5L4Ydq���'��l�q6u��P� ����w�?9rv^f$ax�@�=�N�/ѓ���&F!�f:���I #g�z�b�#�u��|*p�.W$�B�젴aB y�6@[�GXk�� #A3j�yUӖ�8��h�!�5���P��Ė<�� ���^�rV�T�P����2$������W*x'��8�/�N[���`� oi��O}�3�!8V�pP8z:~�4��M�$n��(d�&����Cil��YU	�4���Ġ*+�'p�!�h� P�v��d(\���^�J��x2
��I���]`�M�T�����Ob0Hc��I4�� �i���K.W�@��@(���jAP69l�8 vƕ�ez�GO1� �#��c.N�И}����^	�'�(�5`�]��7E%>#P�F2Q��. #�R�"������0U�,j�,WZ�
h��%菜F�6��T�e4 ��K�j�O���J��{�Ď`�Y1$HE����0+@���� ѱ$�;���z դ���R ɋf�5Cl�$roC'd@ J&����3τ���5B�S����������[�����O���S�LX<[/�5��C`�-�� w�j������p���o��	]�r.�B��ʣ��9j�vK��l�@NC T�{j�e��S��ay�@nKg �ʔ��$*���T������pi����Иhd �ZDڇ��e "��ӓ���q�N �k���M�Ί/��BU�
& �r>Ĕé���Z LB� �M���L9�8~}w�cT��R%(���&�7���$`��	��Ⱦ���Gy\$(O2�(D��@���Ty6K	�R�����&-1�(��@��:Wl �^釽�SP�px.����C� ��P��6�\FtI�`e��䚲��w��C���*\�	"�I���)ȟٿ.�x�B��IS�F��v�t��Ǹ �&p�Zn@���	�8 �=k�mwװą��#`�Ą�+�^������ Կ6m
��T��t-��:0�� �gxw���'V���(�A�=�D�Q���:	���>bǉ�i�9�b�������T@�^(wur=p�'�9�v��eW�1_�~f�H8�&� ��')��24��6��`A�
<�(���rm����� n
��d˖MR�� ����Z9�.L$�E&g�0E\^2�D=�Ep���F��fH&�X� 0
�80���L�!h-�e��Y<��K �~mi��xZ�X0B�  ����M���`��\$���Ph������~u�k $ �2*\%WN/\��DP���x�(����x��̌�:\��M��D,<�h �j�E���t$��O? ^o����M�:Y%X�h <Eov 蓷Ĭ�w����>�j����'߱�������Q��X���9�)� xj	*�H��$������PtF��0Z(W��`x�_�,TB�K+P@��\�����빈 �|>�I�\���l@�i휚ð^�?���� j>��}[}0Qh(���	SzT�����x s;$�R �5�p�D�60Z�O�Ot�XqQ��	1�Vt�mÉ �M�Z����wZ ����t�ͨF���� t����R�%+B�]�N	q@�o��Lw/�)'ˋ�t4�x��C���	Pq�y�� �Z)��+��lI&���C���L��:Aiƃ���9^�%Lkȼ>� ���w���	 ��]a�zc�|�7��������p�*0BR_� �S� �����q�i]�$�%z텐΀����Y�{��>Ǚ�? �T�$��H ������%��&P`a�P���:������j�]����R�Q��H��0UHT
(^�����:�׻ϗ鑂����+�bŒ �'#`}���ˑ���� �2|?��5>W���L�� ��?������{@`�=&�5�9�W$�X	��@PL��0�ށh�` ���d�z!� ��$m��;P�L�����4/k�p茀��+��\�ɏ,$��i�0d<`����Lx�B�	FI�@t#@Q�=�j�����5�([� �������^F;,��~�?��t}�%0� a����X ��j(�9���;G�8 &���
��`(q�}��<�{i�l��؈#�!���\���L� ��A{ZJ����/(ِ|�z��J.�## �wVc�\�I"�>�H*�I��PL<%�n,�РH>�JJ�X��* �ڌe q��-�.;Bᄿ�0��w�@Ԛ��r�8^���Z��`�g_֜�^!л�?^�jT�(���X��@LwJ������ �f���@�z SDT�V͜l#�9�`���[�AX/٧��;�l �g��l�8��cuE��XԣK� ��`��(>���w,�� ��s��j ��Ua���yP� S���6�RK��� �Xw����2��E��i��[�9����Dy� �fJ&?�
�67�ذ��2O�G�WM��X4� ��g;��[Z���Z L��u��i� �pOc.�����'휺�TH?F@l������iOhĴ�<��]���T¬�X(��<�?�u�[�`S)��g}�ϣ�#�`�u�M��N���.�����af���@���R�@
^ќLZ��Bb��_"�`� 2G���$������a�EѬy&o �A}s�U� �������t�	.�e��7���&0���i�a���5��(�?���8���5!��@�	��$�v�@����q� �2�/M�vV)
���� �녬Q�����RNA����- �#����NlЃ�L�` 0M�-����Yϒ��� H�Rء	-��P?���4K����� �9f�T� ��~�RY�t�=� �ly��3 �\�~�H��&��t�{��~�s+K�L��UJ��]��BF� �u4�dx��� �IA[��kr��� !�����Y���Y�O��.X0R� ���1���G�\����� 
�y�-Z� ��fW�팦�m�' �����
<q.3)r������@Hjkf�v�N(�������d`��{�M0
q]T� ���m>lY����F\
�y=���s�&w�Y f�o �m.x�@����҈��#
�ޘ���?��d1������C��uq6����v����@S����g��@��Î�G�1��R�Pq"���0���	�ԑȟ"�y��c�� (��V�ɾ�N��9>�Ro-ca'�	�+I �:=�zNqG"����#+	��7��(���&�Gi����Q�(5�trDdh8�F��1 ��9~ْ.�y2��G �B9�4
@K΍�PY�sf�5Gu�Y�h���9��F�"��9�X��z('��"��j�a���I�&�(��z�H܅^�>G��?�:��.u�jE�Y���o �'�S��������0�S��\e`��ksj�h����@pC�)~/�b�"���~� �[Ǿ���.���� o��*��y2�0!��o 8v�m��]�k���N `���#C$��a��Ϩ 1��[�����J�h��vĤ<T���{;�|�ȸ���o��FZ"� �o�`�cv`���͡@��yI���Ҩ��n��~cO �ڙ�����j�Y��q���y�=!8� .@'C�*�q�T=��I���H(��i�	z� Pن{�0�
8P�=&�dMk���`�[t��	�����0�9}�Z����90�q a�Y�?�.D- �lN���I_f�ȿ�D�U�z���s�(�u`�	�!�;�c�A�S���` �dJL��q��/W��Gt1r��];e>�\�����~�F��d?8�&C.
q�� ��!@��%��Ikt |p٦|�\�(P(����q�b;$9����H7.U��qf�4�0x�a����`1��h����q��D?3�&!�*��~①8�Ap�`��.d�G��������x��F.X���K���qo�� m��k`I��x�b �a?�K�B�\�"�@�ʘA8����#u����Q�a�]�Y�Ȝ#��9|�b����9�|o}�Wl��`�Io;��[ңwU^��.WVt�� �MU�tN9�7^��8Z������6�2X�yO J��q zw� $�(oXb�!Y{4 ��W������C0�{�)k[uP ��s�	*V7�/���)����G�kM���J
@�bQ`��wdq���Ȁ�9{٪� ��9UI�;�
������ Ѳ�l]1Z`�􀏝v!��C���0T~o��2���o�� g�喿���mN�h�q�4@��{L�r3�0�m"���]�yB�Qu��`#��9�ٺ^�Ƚ9g5�w �x"	Ȣ�`(�1(��z��O��bQ ��;s��u- y��*�6|2w�Gl1@����Y�����`-`�Ur���$*)��.W2X�1���uF�"�9�耧��Y�5	��.  ��� /<�&J�*7����.NX������I��8�`�o�������oG�5l�#iI����{�� �Q	x��� k�~9�� �Ld���ɶ�u��b�D$�vp�1Eˎ��������< 9$;G��o7/���P���Y�L��� ��$�����0��,'�|dE@.��|���f6vJ_%0�� M�@�;X�u�7p�@h:Z��_��%j���&V�D �c��~����)���R��
�g�����O~2�X,"� C��}��
��.��&u��d� ��e�Ŭ� ȧ�~A��L�����w~�d�uĤ��#f6H-_G�Ƞu�I��K�̑���b�u�1���̺5E�Ր�r��]��;��yk@Ǡ��w���C�z�YW��� 9?�Nj#������]��D�� �����Q'B��4��ڟvK�0|B�P���s���V֘]�����q��=|1}dȹ`��q7��A�4��� �.�{Bk�X������ �7��{��!p'�M�ל���y)P��j�z-  �5���m>�V8t#b�L@~G2�A���I�sh ��ƺ0����>徤yP@ve� �Z^�ش48� �����I]^�\�xƂ7:	�v��y�W�YJ�ɏ�&)c��_03�� ���?q��d���b%`l9z\�GrPTd�()u2d�7��I�žV| a���Mu�H2L#� ��q��D>2 �~���Q��[L�^�q�~c��
���}����}fp ��/��� �v�FuOH���;OkTH��
���.��G� �����x)!�1�Gk3�-�/��8��@$p�@&��d!u+%�T���G����|�y�k� �	�?90�y�� \F/���0`T�x� &�MC�B�y�T[���d$Iq�,��7'��D��Y1, ��Fz���(�������|Ѷ��r2����Ƕ>�u��hǈ�0jI���e���x��0�;0p� r��f���X�;0�� �����M��G.���{�l����,������E��@a��*Jތ��ʥ���Ћ�q�@�]��\T���	��fҀ�e�������(<��_�,zrWhMc��t`��g�mC� $3=��u����
��Q�o�����n"�TXb�C�[�d�$z�Hn��-�dIb��v$�k.c$���]�����ܔD��h6��-D󀠑�cN�t�$]��#���R7�m.Sqq�y�����w�qޥ<�xb ̩�D;`Ӥ����w�^e0 �Sw���C��Ц�J�A��.�G`ԑ
Ⱦ�H��[A��1�Q���k�,��%� q.6b|R��D@`�*�?���u���Lyl�Fע���V�b 8ɵR��k�a8�-�T��{�M*�(	B=��R)>V���	��� �q�\jxf` ��y���Sތ�&���� u��ʗ�S ��NC�O����K{�E@F7�`��d�Č>/��J�4 e�Q�/�b��5�_�P�Ĳ�a��2� ,, �����hέ���.)�yn T_^���+i�ްXȢW�7��F�!H��1���u�38���o|�`�w�� �G���x�,�FP�Y����A�P��j0��u�Q��m���i}�S�%�����̃� �����T�P���o8]a@�2���@�n�Yb#�	`�s|[��0�o����������0�k�dܽ ��DB�MR�;-���}	o���� օo�Gr����,������-k����:�#>�0|�0([K(�MD`�8���z�4��+;Y���4�=� ����꜅�� ��M���]�<jQ�����Þሚ�a^�`B����!�� �ȕ��y��
��q����{o��z�D��oL���yT�9
�G�.|\F@ �>�{K搬$�~-$�A��~�}��c�Bm��P��(�u��0��o^�ؤR� ��\���͔�|o��bC�" τo}ٕ30k���p� ��(�lŰ�N�u	���ь�����(0�#���Ĥ茎�@u��^�L�T Y$T�J�%�zH8�� �"�cx�I��Ѷ�4����D�ސ�ˊ��1�+.D �\�P�X @�5�	i� ]Z��O�.�?K� Br���]u� ��n������(�K@��0� ]<v,R��t�')  9�]���=��W�� �.��s@2�wcN�ϐ����]S7�r�+@�=�����P�J��p�?a��O����\���11�1�惘����8� #?]��K����(���v �9��
>�K�6F$�Y��XpW�3P/Y� !q�X u�MHS� ]��.5O��0�P��b���q�����:�xW�|�)�/O� (f��#t� �>��ux
�Jv܄+��S�^�����˵��|�]������9��%g/B����(�L@�]!vDb*$:�e����T2�嘖Ed�#`y���7�%���.� @�z�)ܠ�{�lL0�>*������-���D ��XfW���@o�X4�E��w��9�H��-z�*ҷ4���Φz<,M F�hb�7[8�f:1 ֢��F���ə]f8@���4;�S� �M��`���<3�d�U��`�1��'� �f6��#�d��=n]����| ����ᰣw �Mf����8�eW������Anp�� ��~m%�HE /����+=�h�d�0(�S�� ���q��8��(��9�t�%�g���>�0�FJ#�g���� �?�� ݮ{X/�;�$D|
S=�|F�:4�糸�8�?L`X�_����+Vš��Uv,c�<�0j��q2�Р�+\ V���;�t !"��/+�3��% !�*��ǫ�{���q	������i����F$E� �5;�[3�L�4��A�̂�wCk�DD��TYz� �q����J��MEb�`�y�'&0�x�P$ܛ� ��,;N��)&Ö��5/ #����"�c��j1>���$g\ڥ�����L�
-dN��� q}��!>��$�L	$��À��> )za��UJ�`ȸQ�Bo���C��r�O�P���]&v�b$ ��]A ��d� >9�\^�VPǠx�F�d��K��<�q���b�T�Ĳ�
� ��K	�h0��� �@g耘��y'
Zn`׊9���x2dA@؁`�i��z t3Z߽���x�΄R���5�x��c�ζ���:&`�g�a0���)��"��2T���e
��<@P�=:��X��s�E$�1Lٶ�Q��S6����r���(���2A��c���L�|#= ��9�:�M�0����qo�� ��sw�����8�V�+7�Ki�j���,�"��)%�Fv�jA��b�� p'���`�o���Ȕ} x���)���	��2w X�ݙp��� 1|�C~ݤ�9�����@�bp^| �v���3���=W��P�N��	�o���m�:�#L8�<��$�(�#vt8 ���] �ޓ��W� 6J��1NQv�{�P�W��H)~�@3���0���.8� �δ<P�%����� `��R����_�g�-(�k� 6G���Na��o�h�`W�8�8Jx\F% upЄ��p4^AhF�w+�e�N�#ë��O���]�&)D� ��0\�>��]�P쫳(Z@���2ث�Oj<"�(��;��������Ƒ���]%v�q��] �P*q�4>�\S��LȨ��̆���h��] vF�") ��]5�_`��N"B,Y�����!�� ��� �,=nW2��`u>�t��S�n ���� ������?�T&�I��.��g���x�G�5$�(@#����OA`�&�s ��ԙ]�-��֦Џ�q��NI'�%����R�wqR���ؑ$���M�i aD�*,�Z�8t2�"��0�]"v<0���]�&T��R�οԊ�Q�ͼf<�^*o�� R+ 9�p>vc�H�x���9� {	�����
 W�rYF��P/�O���������*��}o�H�3���gbCt��(���0CJ ���3�U1β�GT�,B�(�X��#H3d�q�����)�0������Dd�J���̈́RP	�b5�8��c�y�5Cx!j��=d�(��XdWF�"�uX�ס�R��@]�r�� ���U3ҵ,#���;0���G�w��inE��8�'�$=ٲ� ;e��� I\���+	>0��΀����bq�����RF�#9����=�7O4D�����\
D �i3�Ľ��LOPW%��+0�XgW���`' ��B$
w��XE��ל4�0� �a�$���0��!6  ��L���z�
��F�� ��� ��v_E) L���[��xy)��� 8&(X�<�K+�#�;���*���(W�
��d��V.�k������� �`R�3�{ �i�r���>�P�d��h�D� �v�:�6
�cm��RqY�# ��"4���EP=B�ς�w+{�S��Z$����ٴr�
dQ�A?��0p���h��h�{IT4 �F)J�� Ak1��+!� ���/��4�E�X��qL�9<�m�Q4s�)�CY,P[x��y'<F^��.,@-��ဘ�c�+Ƈ,�j���@g��ـ�,76)�4�XqW��&j� ��~�y�*���^>�����y�P�0$/~��n ��r�Fp��9��Y4P��� �K�Ѯ"͑������'�˪��W���@�A?u�(�� 5B2F�>��D?�&��ϲ��.�# �	V��c�Z�	��d���Z�N��:�n	��$��(��hݩ�& ��_J8��2�|L*��XrW
b�%k��pw"E���/0閐�?A<ǀ��;´+(g���bh�8 �u7��� S����.F\��U����w�M�%�u�؏ah��I�`D�� ���j�L��\��)~0�S��- *e)W��nX�� x��"зd������(00`3�Ơʕ*T�MK�a�6��CpY`��ӀhUw�L9�P5y�7;���S������ 5��U��Ԗ�\F#��`��I���	�'�� l�n��=�F�]�tF��
W��9<zc`|���[o�����O �qb�������d(
��cB�T��'�q��p�%OҀ�Cy����c��B�� PD)+<
 p�����h�>6H%��'q`�- i[AV%ͷE��_�GٜJ����-w�\�⇢��3%����b�/9�y�9��0����̐�C�z��B���@�� �@o��B���J�� �3)�O�t�%��$��0�nX�A�����C]s��L����$�A�1�yf���'N�PGtO���}��I
7b��(9JI�)��|b'� س���߀!8E
H����wh�A@d	ˉ*�hW�&(������A�j�up"���0��?	s�۶D)���� 9F��cKv��ڶ��(�� ��~�V�'b����(�p�U��t���0�*0�=ܳB
��0����:4#"y.䬄���r�	����X��Z9�׭�G $K|u~wq	V�� r)�.�pM(�n#f �����Jv�K��<���0�H c/X��'�0�����Y����0 �Ff�~�UJ.��c^ߘ0p�00���-���#)`��A �����8�����F���]b�L�\tF����5��!,���v���}�O> #�p��7���  ��D�c���JlQ�y��	��� + L����.�0c�:n� &��@Z�-����AnpxĠ�;]݁g��H���C(P�{���. �oT8�C�* ���-5� ����eU��V�������3�xL��P"�`4 ��\e�?7ϰ�=5�	�t~�QD���hhͿX�+Y� �z&p	S�2���XV�\F' �ڿ�5MA�h��09w,�6���O
�5���� ���EHL.�9�@��	!o�p$�1hm�� C��Y��;#@W����N I�1�+F����l`��4�;:5�D��� D#Y.j�@&{��}^�hy�f o�����/�2,N�j��+����ڋ���qW/@� zQ=��v[/J�����sD�'0��Ss桄�"����1� \w-�� ������܁��]�>/�n�H�NL=JfΩ�(���b�hҩ,^]c���0^-�@�L���@6S�X&g ��>N��U���6�@�/H
 t�w�7B�<��0�g�P �JZw2�}�9�6�� �y�\T9:7E��*5��x�$0x���౫�	��O 0��/$ׄ�j�KB�y���~���`!��̯�!'UXog? RK���;$��l�y�6е7� a!�<h�0L�i89k)6�B��~��lL|F� �89���	F]vE���`%��%ٱ!@��k*�] �W���(Tz�h� �_�dٿ���)$y"�s���pB聇d%`͏| CŰ��z[$����]���u��f�� s�/P[J�CP�`<�$���q��| �{#ٸ31�ywS['� �C��B�:h#$V� �q"�h~�CB��֕�G'0/4恋3r��ƴZ�/�#) ��9����l�'ע�]p�e��� =�#)$w�pA��S�F��~� g���>y��{��+�ߟ�%�N�� Li�W���v�<�H� ��%��k#�ۋX�p\x�-�ls�X�&� B�TA��':A�)��p�nm��H�ܼL�-"�5jd��dD'`W�s��f$$�� �������5�hD�w[O�K���9� ������'�쀷�x�����'e�������@��1}zt/9��I��c�*���7� RA�O�lNy��� uC7�ZK:�##�S� 7>[�����t0\�1p�����
�ٹ��D�'�B��8^�	���đ�q��*�f�]>\t,��	�L�(`�vF��Ԡ�4]���B��D+ˬ������cƓw6��!S�� �1�-`*����ԟ�')o��2�a(�� �(ZK�D֛��F� 	�V<a!������@B��ľ?/L�o� ���qX�J���V2�z�!��ϓԀ�y���Ш��6P��������k��Лs��&0qf� 䆅��Ay�$9{HX1\G��r�r8K6˴����]�q�+�£If7�y��w�������%��<��q0��`�&s� κ�:�����+����(0�+j�2�7U��..�yC)>H��쿪���9�(��=R��y"��B�H@g6�[{� �ЕY�/s��< ��y��%g��-�1Z�a���#�\@�|)�)L���S[�����W���jX�P �1DH�ƛ��p6�w�p�0>N8 !=����S�>tD>6̝8�Z.l#) O�\���e?�r8]~��������3�{�"r��c?H�8w�J� 0,b� ]�� ���3H��)d\ ��l�7G�hz�C%L��3�l7�M+���Ŕ� >�)�B�r 2�pf�;��?�9$%, �����.�,i��PAE �"F
B�b0x�����[/P�,�X���� 0E���`�Q�_z3�`��)�n�;� R���
����;uj�!��L 1����o 2F�<'9Y�Hn��J �˸�#ãаD9�L�)ٮ�=�β�4+��;��U�4d)`?��([��+�!(���1��������4��D�ہ�W1m$J� k������,�h��s15q Q\�ұX��r�����n� �_�6���[&�XTzE� T�u�w/�~�`�7e��`ʭ��l��*	ٷ��.� 9i3 0��v�c �Y��$q��p���)��!�ܼM��I�ճ�������l���(�}�j/{��XkV-Ss�>� �/��������b�Zx��:@�����	KV��JP<s!'�>+0[�X��ۇ��Fb*�u��%�p�~ H]��*�J0��ac��`D"`4$�J��I �f)h�^>��p��	O��p/3j� ��hbĈ�NW��U��8(]��b�vS��L����`��>�c����iIxQ{�`��^��a�:�DP��z��/:�#� S��~��j�˻#��ǌ%	�����5XX:��<�H�U8?�0��>o� �SnX�3޴�j$\�� ����C�%䶡NȠܱ� �E���|(��,0���tG�>Zܬdޅ� h��g rF-�sB�� �7��#'�'�!���C�x%BRДJ@�4v-[��t�E��>#�=�D!~�$�	r�T@����@��(X��Q% �S��z�I�����(� P�����8�Z=�pG�67Q��� u���`�]��ǴA�C9�pO>�#� ��C�vp}e��lQ���� q95�Q2�.<�$�4��J2�4-6���ǀ�H��\=JPr�+p:E �y@�h���K?�Y�\�x��F�Lp "� ?�I/�vc��h��<"
S�ie���`�|jU�vXK�h f�u'�x`G��@�]�z��_��� ��R{$��`�0n�ctz�<&,K�H���_�� �b���<�}��!H���|=3Ҍ?�. ηA4���`7��91H
��~ �MQVC�  ����k�ø1���XxAr�jP� hm[�d̆�\�#!�_ mD%�� \��ޱ��� �v7mq��� ��w��a NG��4��b9�Ł��_�@�&:ڥT�)c�wI�Q���V!v�x�����.�TX>N8��Ҁ��W�
'�����gլ�A�e0F����E%$֠䃥[��42y���0gm`�l��zbm�L&�@ņ�o�3
��fXGd�v'����\�O�:*@@ٳ$n� ���X�	s�\�m"Z�\1$�ħ ���-�Um6���� ��ϣ��$�0&3�}ï' ����sJ�������m�w� �?�%�@>��f(�! �7ݒp�Og�`��N \�ix��m��we�!* p���oW�<3���(  ���_�� =I|B�h��WVz��0��E��C���)M�2��l1>�$�F8"� �6� �sT��h)�L�-���[#2.fJ��_�"�� 1Q��a��:)7D�F��2�!a!7���S)Uy��e�~ ��4t5`�8�̧�S�K�`�!ŧ=��녀�\�z�l64 �n�+�� k�w��V�0��QS1�c'0�#�6ͧDS�b� Ƨ ǩ�\��CH�<���_ީ �����ȅ8j���D�S:��<E��l){���/0΄a{����ƀ���tϯ��M����0��7ԧu#S�� ǧ���p�yD� �g��U�`"�E	����!��̀Q*���΂1h��݀!�m�	}�?*[��
���A��zn��Q�˧rS��D�
�d Qlu�Sfeh���j)������E�\����S� ��iL���H(
CW����9���;�ҧySC���	�� �	��oSڔ��0\{QԀ��Do�Gu� U7p�0��y�;j�@H�$2�tÀ"7=��D3Z`Xlv�� ���Hy�U4p�+{�K1�D�!�<���(�Y=D|D�0���MY���kc=�#�0� �5�oOKy�s� ye��&�!�\��1�hrz�d����(7C�>�Q` �����!����*��)Pz��i�x{�}�y���z���t#��#7>�6�b6@HmL�ߋ�5 �߄O=��� ��
u�P��j�z<"�(����4ݰ*��aVJ
����oOL�t��mnb� &l�_Y��Qj�CB��0$7?��1�\7v;WC����L�(�H<Xm�3��+ �ٻ�y��$Ȁ'7B�6�(�_7x$��A�\�� n��%�5��S|mfb�� %k�hD�	��K���ր>�#����� �Q���j姈�4`����r�&! ��t!
�(���LjZmD������$�����T�D虫��O١��q�m��;�~�,��� y}PE)J�����|xPO�q� {M4�[�
J��D�`�25i�X �y�{ �4l�����k �<yZ��Ip�B�(�X�D�� :�}����\Nx���� L�k�|���o�c�}w�N��d�`�N3 2����7y��0���CD;k��� �	ctlr���g��!�m��<l� ��6S	� �@�w@ �G��D��{�`[����mFa�M�[�  A��!"��i/�|X�؉C@4�jJ��:�#0 O�ڣ*���p�`�1����tTW5�(	 !�����mN�,P+ q��]�\�� Cp�N��|����&҄8��������Ja/�#�r���D}Ͳ8D���%7@�L&��]7 �W���;	j��{��)C_H�\FE��0r��m^�$j�?}K ���2�q��f��q$�9`Чw!S��ɧ� 0����j&�)M��q��'ـ,t�[Ӝ� Unf=�r�5/P#�0	�7���fB3<'	����a�y�)x^F3�L������,B[z U)2@�4D��Ȉ� r��kcv�M�)Pt�)ҕ+��L>�B"J�\e�W�/�#3 ^�q@~ *l��+$����YU:`#5 ��Z�.�H��0,!ˡ ��A���nⅮ���XV�%g��T���0	2���)H��D�cZ��s�-Qp:d�kxS��X� ���P|9q��U1]���'�h �o� a���D��������juUgF�DO�0u��mv,(�'荭_aH�E��K�Ȏ����2%x���Ĩ-�'���u��p�A����7)HL��8���A�8m��Uo�V^y�g����d6��HZ��3��	
�R"(�1���c���0�$P�r�I�l�!֬�\F� B@��)#��;����ތQ5��J���������3`�50�P�;L�@����7ё `j��	�6)W,�C����q�Z��͞��(�0�<���i��rm���\mx ��ז�060]�8?�<�M�)���^ՏY�������Q�d�!�K,}���*��0���g=n %� �.���U����R�E� ���i��p ~&jD��;e����|N �`7�wY�	�|���\xp(��8�2X���9��y��i���{�� KJ~�f�X? ��0��=~�yl��6n���h��@:lBB8�61��� ���G�u��0���8��� mc�}K��')U��ހ��&���tF2�y�c8��:jC�TP�A��4� �uɩo���2pX� ��I���qKB�Խ����U�y��*�P�docA�'�P�D�� 9ݛnT�� s�7���)D����`��xH슌�,�Lu������ n|����ә�Ј�����S�-tM�`�{��,ߗd�u'�� P�oBp�w~�0��a���v���$������GjK�/�#.Z��
 ��+���A�r 1q(�����	k�d�Ǽd5`=��P���o�c���0�;�	k�f�CW2���^^�#�������lr�J�X���g [�. �L��ʪD�Rj��ysm�\� U��;=�����M"��/�B�h��K:~��q��8P2�x��a�)���
�t��3��(9�5�9� ���GQ��1�*���:�h�i��JlYя"$�� �Kڧsz%��O�@zV��&	���Oqd�]�A�}�~��5� �'iWb���m�#u��\LQ�tC�)�` �;�9
�J�瞒������g"��`ڋ}�_��� U6+sj,k�؅�t'�A��wK a7N�}D)�LEM՗pϬ!y�5x @�gP�U&/���(8F~jIy�$P�ze�Kʏ�����[�%��i����������{��0K������#1h���Fͨ��7( n�P<��&|�"�N/(~� g"ߏ?�J٭+�T���62`O�� �����0O�
,�`��L����;x��W-�����0T)>L�PJ��j��p�X@��� i��5%�T!��)�s�g'�ӓ�uΜ��@���p  9���� �!f�:TZ�4��숌��|��� v�^w�
������ZU�L�	��w� ;��)�jn%��@���7�*9 7�e ��8gvW��y�	N�O�����%�/�)�mĸ� � p-D�D.��/@�0�\�` ������QICgu�Ҟ G��/`4�U9)
H�o����/6�8�����hOy� eK���t�����W����KZ�eS)�C�wj��0m���x%T�<7����.�#� �uDe�	KB�����Jӈ (v�#)����JP���l�;�Q�q��&�g� Y�k*��`�q(��]w�${� �I�����	"�3*.0Ǡ�Kg��|4��~��aoH9���^�A`03�� \O�5�;�ۻ���HGp��{ld��@�����r}	 ��0k�)W�H���� E��m�/�X�0>��<C�K���u@���-�h����i[�3�� �KJ�ג�����������x�t*\� 1Iܔ>��n�OUQ���o��x�)p	F`�pq`э�~� |X1ؙ�6*]��|���T�M� ���]F�� �?�����>&��ptF.��g�ذ������Bc�A�T ;njȢ�d:���L�0iL��q'�1���JI��f� (�w��m�b� )o�?Yd/�$��Z]����d�R t�S�TU4O��\F�;U� ӻJٓ�eו%d����Bl��00�Ѻڢ���j�?�|��o�{���sQ�+n� :�ŏQ��=�-�F0C_�K�����ӄ`ºh <X)Z���.W���2߀Uf�D+I &x�WZbk��1��A�G�U��(�e��(���0E�0\�݁W}9��"Ao�z�*A<×�kDp��@ �<0�%�c� h���1�"�NBnt >�N���S�5@�g�8|F�>�܏�#��G��� �k���8 ₛ12�ݡ�^�	��H��r0`D4#�9D �t�r�Y�UJ5�������~,��'a�3
��h�pD���`|z���1`P�oH�''j@E#sO�<X\���� �Y�Oi�$����*2� t��E�Η-�C�HJ�����ol �O�5��$�� :(W�X�	}g��Et�`�ܣ	5��qR�jSx)P�1٣��h�_�X�؁�	R/������>�i�0\��� ���G���(dx��oϯ{
�GO@����]��dG� �g�[�8Z5���.�r����X\Sݢ�����T�`�M;��Bb��d�UJ�����t��8 J�/p��Q��m��%�SmU����Ҽu Cg���|�ԑ��y��Uk������o�)V0ipW�N��x�=V$����I|���Y�� I�g��[�|'�H=H�(K������s�Y~h��J��ˇH�	v��$���Z�"%��Aknʌ�bKE�3���Ytl�w a02�����t�����o{\tL"�,��8O���������`��xϓZ,\:P#0c�mi8	#_Y��-�h'�HH@����Fp�8d�	�������\�f��L���$��Umxj����]�e�Q��X!/Ke���`�
� ����3 �(uq˰��t�O����.k$ Y�g���v����>j<ݹqj`|.!�CV	+�g㩌�t���������B�y �-���J��bd��|F1 �jZK�Y�o�������)$T����K=��d���O.��O!ȂqkWز� ݊��BbÞ�'�� ��'L-@U1�T�NK���d`�����>5���)џ� y�އ�� �Q=�C)�Xj$��ڸ�����,5�?����J��pmr��>��:|#� �Ӈ;$�K���LXE
�i"N�)P����,���8z������\�a���C�1zJ �,���M��etY�4
Vp���0Y=���O��H�	�A�ߥ�:#�]ҳz�Ȣ�-������ &t�7��  �zm�c}���4�T��0��,�TLy@�e�k<p~�la�Sex(�����$���3�R���XՀN�*�rd�
�O���y��� ��E�Kk陠���� ^=��<2 ��|ː� #�^x� �������(����ќ�.�L؇� ��Y�yKC�3��0N�<���Ji��b��Sa�?/;�#��N(��p3@yS'�����]�Ŕ��`���_��(�O` ��Uw �8�+�W	�S�V kM�D�4��� E�O�H�p&~��	{(_���\�1�x�v�(ļ���z�p�T�o>7<�c��Ќ�ueg��'����N2 �[5�UknZ�HȊ�^�UnO����0������T�/� A��j�|��t�& Z/��N�G	���=	T���t��ɉ�����@��CT��Zɔ��ׅ��5ȼlJ;���]��\�� �����"�9мLk��ѤJ���r�GY�$:�#��#~������zU1KF��#�+�p�m�@�
}�@�E[`��|F	ЧkA��z_es��*�4���i�bV�hEm �c��U2P�$�0<gT�	R�	��8��*�`ϋ X[ԿM1�_-�} �@�7���C�Q�=� g�q�� ���"��#� �] �s��3��mt�B��*"�%��(��{�:�0�<� �)\�� �G�y��[`���0�����)R�<����~�����qt��YF�)�U�����|���g��|�Q�X P$9	4�E{��,O��Һ����\�W�xKyy�� A������$*1��Ej0���x�����.m�� �?-z0��Q7�q� {�=MY]$,����$�xd?Q���ɣ_��$WV�z������`x�Ddv����|-�dˠ��5�L��ߌs�=�yia��<M����e �3@�K�q��j�@c;S8����_��?������>�m��Enճz)P(�����G���݄�#W�D�YU��I�I�f�
�_W9r�0?���,v�_�k��	�I������K��Tۘ�w�0�Tҭ�A����`U��q�Y�m�q�R �אP�E�`C1 	��#
�ťςk�
P��y�0	���R���A���� ������F��'��{Hr �M�#_�	�7X�j�ׇ$���"�L^F� �E�%���",�m���pM-5嗌�F �ǣ{19P�� "�03��ȼ������#��8t��$|F �������L���'�m<�B����٥!�P���Ā�pOJǦ"?�g�h\� 0�ͪY/�k� �_L%%�\hX�'�t�4�D���~plo�U�����t�磝�l�;j'_  ��� �(�����J��(�0� �'��i|�/�)O�QT�' �Rȣۑ/����Nrɸ~0������y� �G��U��*�:T#3� ԧ��U)K�8��<� >e{=� /��2�K,�bL����"�2� ��aS�K[@��N���n��B�0M{p'G��X���N��J��*���mu˶�F�TK����S���� �b����I��KP�H ��H(���J ���ϰC;�ٽu�W�8y���#�%*�0Q��C	S<8��o�N; p�F�u� ����{,�*�o��� �e�Q�7AU5�-�é�*` ��8��O���޲��?��
�Cw���_; ��KRnz�H��/�e�6����������P�z�wyRz^|1n� ZX���u�8Nj`f���`+f�P
`��=ha���-�g�#�	+��TP}�^$�.�#�4֤��2�!`�Ze 8ݿo���z�aj����`�L/9%�@��c?��"d�~p� ��T>���B���#���^f��9��mv��}�����b�����qx.f�e�6������	_�QIO��D�Tj͂���}>vI�n��Nc�@G��ak�y%��!,M���]�6I����� S�Th�Z��7lO���'��D`��� \Ī�	��ν��-�1-ǅFA��{�;�� m�����V�O��d֔)�YYU���u�����/��Z�f���
�0Y( "-�ς���#��\�=tF �gT3f�����%J��Ч/��]	���S�����F,���J�a�\�MQ�tm�����>���^PR�"�-�'��B�7Ϟ� �����gHy�"�:�k.�M�`��o���!� �ƻV�k��	�8��p��WߩA�q��n�>y�_ j)@���+� :�x���R�T�����tS�� �$^��o�=ゑ��l� �:���G� }����f��`	�YՀ&�a+��Ù"���I ���XV��Pʄq	�Z� ���s�t� ,��笽_�soP��3e�z���I�����z��&�^�X�J^�:�# p^��r-q}�S�����FbH�]���˨��@�g��jH����$��,a� �=���P��H��HV���"U
�a>Ad$�<�$�vG��{��� 7U��m �ub_��{��Ӛ藔�'D#�Q�{��ꪃ� �63)�a
�� T o��V!�y- <���)⩒�H�����g����=�|61C�m��^��o%��X����*����>����v� !�1G�)�&�f�i�C�g���G������͕6�{ .���;D#6>���2a`��r��q;��Bf�[	,F�o�b���[�5�.����\�U�k���_-[�L���[��
�����+���=4�@�(
=���* ��WETM�S���3�1�IK0t��z�� R_�ir~r��~အxۆ�_ ��:�~ǅJM �}��UY�7���{%ytl���9�p���y���Ku�)�vߣ��"�Xݽ���>�֯�
�;�f��%��),l��x��d���~%	�H$[ ~sTo]%�
*�ċ��y�A{���� O�镪�%��n�`��������ѽ9�'�P [��{�E�� ��MI��-1fa��D`�dk/G�ՠ��}� ����r9!��� �u�^�y�q��:���?m�wJ�<)�Tў`���B����)7�׳�y�� *i$�4�}!��X�◻�Ҟ��Ǎ�ͤ��]�:&G�da��TVP��AF	�����&�[/�8�0h8:T�^JM���ީJ�CQ

�I�y��A +��""e�%�뤢j �r)$�F� �w��ō+�΋[�2�N�����X�S�7!��&��`��Т�	9������_4A�y%����D/)	շ����N�XY� 1���at�$�Z��̀��H` ��af�A[���$�[� /a�>�����s1��y���o���W�g��Sb/�5�QA~���v :R��a�j��7f^�?� q�B����p��)e����)!5�aJ-	��&G/�k�� ?����%��G��/#&�#֋�Y��kd�=1֖~��S5�r��5PN� �T��3�}�'	�H��v9U�?��Bk� �G̹b�Q�����������xMf�F�����=B�L!ѾB��I�6"��� ;��_��=��� �1�XP�� �Q���v��ǅ[�׵:��"��3�c�t�=�On8j� i_�ђQ�JED���%X�¿:Q �"v�k�a8��_>�# �t����,+�!��*��`p7�A��)�� �9i&�fܽ�vC8_�j7<8���P��������H���L�0$��p���i�5[dp�e���Tr �$HP�m13Y�H�[��nf�ib�*-"ql�3̼���i:��5��.���2�A�i�7L Xjq���p�
m[� �ǜG ��_ oi 7�dƒ������^�@�Ű�$� VΡ~y�fp��3��#��K�nK �u��_	�)��1-&��^i
3��,���L%��*�1&��/�5U��[�C������ �{��Ro�\@���D��K;�`H�U,�~��,�e� �0P�U��_Y�#�1�a$�t#�`!��3 zD����a��7�`�����]UE�y^����*ل(`�Td��1ma�q#��0FU�z���3����{~p�Ef�r���[��ֽ%@�f��&�`?���1�EV�C�)؋{v �
��D���Y�-Kn'�	�r�����Y-u���N�3�������򡉝�����=o��~1�)��_�/ɕ�0�dPN5Kz� �OoTK[H���$wh;� =|�(:}����Yt������vX��lR=� ǝ����,%Dc��$��+	��	3��"ڨ/��0(�k9|7����q\F�j�'6���q�fu� 2`�&�?Ha��8���� �Q�6+�)�.�x@��$Ȋ��,g��D ��8�/*J�m�\�^Y*58;�[����a�Cflˍ�q )��dm��4���"B��qhE���l %�Cl�D�x�Pa��p`G|sr]��S��fLY��Nx�'2��!�s�s�������b:{#ku��Ƽ��tI�� �,����� �.jw^��Mӆo �6���Q�����`^���U�k!��M(`�CGRP�ҤQ�"�+��@ͻ���/6��`eI�au0�/�1${ٴ�U�����f`���Ҭ��
C9��5EE�Wo*A�M��s�-g��b �"���~�q� �;�A�pmܓ��np=�.'��m�C��mOK���Ε�Qm3�k���|���� s2p���h���4�@�f���a)鞢������=�S0��b��}f4#����k�!�m�ah_������O��E��k�t��+� T5R&fY��U̾������ 䑾@8� ,�������[�p�%l��~���5D. 6�E) u��@���N��_��:�d���|�B8����� [���T%�D��bs:�# /��_�������ӷ�	�a�^�i��k�W ��TJ���x�l��$�W�ܬj�t���q������o;�#��?4���%������ ��a�W ����>FIP_��%j�HDa3��;�	������ެ$u<�P��|�I���r�p�]�@y�`x��,���a�my�1	2	f��Ϛ1����T�a%�
 �fx�j+�� 'kѷr vC^%������l��]��_�s�q_3n�U����h�	j�� �*\1�ƭ ������[f�ߏPѾ ;����� ����,�V� �)��{P[�%����Ho�t�z,��AjA i3S .��`�|�� � a�����P&WfS�,11$���*nD no�AN���O�|��s�����C^[͗v��F}��Z�j�Ӊs�W�%NǥV��I�����G$u�N���`_��O�0S9�z�,�p�q �Z����1��ǄA�ȉ�y,�N$�����0�qZɐ�J���E(�œ�@�-�8%+�d� SH[���� ����I�3�+���� ̀�K�{�S����0CuA#0���
4��@;PА�(��E�H���g�'�NN`1�%��+�%f�]�����`e�������p��d���;j��d���>�Y#���������هs#��mG%
C�ߢ�7�	��m��J�l�G�
 ����
�y+��Q.<-�MQ���;%��U�e M���#����W��-��3�g�n�� �u�)�p	�^�[-!�k�>v���b��_���w�q� '��7ʉaT'ĝ��H�]"�F` ���4�P�r���J��X�Y"�_7o����;�׸`�������a��g`�8��-�KI$ �5�L-�ጙ0 A���1�Yr��LE��n�)��E����}1��\���/g��S �D���;1.j��)�.p�& Y��6��Ɯ%V�'X�sA�=�H`M"XW��-_��c�����F�<rZ�XW��Գ��8�d�[A����K˕%���	Q�r���3�A��+����nh�� �u�rJ�<���,	1������a�l�܃���I�
�]��j�μ� H��7��>�;:V��@�_h�{4$�{��p��T����}8�Cx��
���	F�[��)�7�Y�a�~�W7\L��`��S�ّ�_ A�Ź�2��e��Q���704�����M�5����D�~3�u!���3d�(�U�rfa����� �%����`V� ���q ����g�X	_a�7���-��)?7P�����SA,�z ���R���7Y!E3�$�TG߉F�@fd�v-� DtVpz�`�����Za&[�('� 4d$���0Ơ$9��?��''E_F��{��@0���������!%��![�a�*˾QY{��a@��$���"�mĉ����hj#�j��Q%�%d��.�Սj
s��r�����3��6�P��N=ng#a��_��1��Qǅc�k5m���*��aY[tD��������_ �P�� '.��,!�,��,'O>@r�����!�3Uz�P0Da���g�L�XZ��66�ds�,fP)(!�X�W�����K�4[fF0#�	����}i�e��s�9�γ�_���k�dmj�x9(�&��O-̫��C0[u�J�}A��` ����vQ�����5����`��� �K�a/�ր�S���Q��,K[���jl ���׿�K��Ƌ���J�� �5��Ԅ�PV�4���,/�"��M�-!�P����ч)Н������H�Ҧ��_o~-?Ȃ9i.	��Ѹ	]���-MkΉ��* ��̓Y1�Q/{/�`���a茖b9�¤��H�Ϻ�b�k��F�����P ��9�B���%	ɖ�Uͱz�¸2��y��%G�+nY�x�ҭָ��ue�>��BU�. ���� ��ȝe�'Z|�y�n|m�?	���v Nr�D@]�s�%���a�5O)"M�]��%�2y_)��lL�I"�kDc�-b\�}��c�%��	�����yP|q�a�>���	8Y	��{��C hU;�a�	�(3��0[�DA�U���%!t���]7` ��f�r'��\���o���u	��	^
�[��O��K�P�v$q��.�*���{�.=��H[��@�������q�qJ�D�.`�:z�����)���P�'��J�BH� �=�����T��(����n�\_j�	�qeks�Q8K�����!�zѝ���=M{[���MS��>K_�I8x[�1��f@&j_�`��<6�'1��\q`�K@���w8�" ���#�Ӌ�a(���M��^��u.���P�Dz�U:J��w�	s[BbqT�D~ �!QhE��O���_�ɖ1�� WxK߄[���� `ͱ��vLG�0��K.�^P�KE�:�]7� ���`u��6��L�P� �^����=K�32�9���/��p�y� �*�p	�U��%�q�7��YA$.06�5�L��)���1��-	�1���+ȟZ��ѐV��\�W��T1����	�q�\I޾$	p�:j��eM1���4)���]8���	�ԣp�=j�������� /애a�ϑ��M�l.a,�M�"?2�]�À�p��'��� �l�dڡ���	P滜qZ,��o�	f���>����+����}���>a%'@O51��%����[�iҠ� ����)Q��S ��w�ON�K��-5�� ��/`1�H-̓`Na4 �x� .t����O3��	Y$Zt�<Q�M��f�y�r(�#�e,���.O�Z�P�5׬����1�.4��0�`�y�i獂g$�V�P��OAE�g�%�b0���
,B�^&b��\ Q{�s��`V�:%WTZ�J�%���g�V�$A�O��V�f�%����R��/�W~���Ev�<��8J�#R��f���,��.ޮ��=��M�$[��@ސ�vZ�'%��hoP.�?!aY۱���ŐS��AJ�,C^tD�-�	j�hY���������g. E����+n��fVvm���s�o� �����9�e�П@�+<��F��������	_[��5��H*`�9�v$��E�'�P�Y-�<$��I�������0�5'�%F����F��	�@PV�O�ڄ�`� r��8�)��퓾R�KS�p�Y yGx��J��Z�Q	hM�2z�$�z�� *B�Ilt�ά%� ����P�v;FZ�]�vI� �����H�\��p���@�i�a6P��M�BQ+=.j'�X�QW�&SXx_{q��D"�.��͎�B����v:	P%�g#\�H+���y���u,Y\�m
���U�:�ҷz#Ra�ץZxQ�K�#��`���2g|i�* �f\-7X�+|1)�[*5��&�' V��ǁARZN���0�T+i�K?�_�ݤ8 z��0}����]� M�:n[_�����)�ݖj ��3ePS[d�tF"N�T��G?HQ�����=��ځ ��m���8��`�	A�5;aҞK���,#��p�R;	�_Q˥�B�������|Fz�:���P=@��T�1�Y��&�J{���r��ቍ)T��TX��S��;����]�
�NC6�-Z�3b>���	�1w�2gtn m�W�����[+t,�j� 'my�V]l�K���W`-a[��4�EʵT�U8�J�&� �ϣ�y�E%�Re01[�p����W=���P�Ca�g5;�u�ٕ��8pA;�H �z%��f��Ru6(Q� � J_�1�J�''�o�`N]��c�OY���)v���J�X��B�T5-sTpv���	Q`Q� 8�=]��(�)@0�r	�
���T	a_Yvk�� �Ef���V�qoH�J�����q
�e������K��'��Vjb��dP`�@l�#� <3��m8��o�>g8�Y�ǩvK�Y���@*z�� wikJ�j�M5��A��?T�N&v�1֟=�ވ �#q�i��k�+l��KH��p!E������cd%L���`��-�Yl/͂��%.${�����ND� '���V��b0��m���%Հߴ��ױt9�$Ѭ=�"�U�i�_m��w��)�I-�xJj
��D><1��v�d5�S�OP�Jz<g��������U"�����>@/�푛�~EZ�,o�#*��J�������	0'e���*�Y�Y[���H���	�Q̉���@���w�2���Q[a��'�4�j��U�;X�V��ԇ`�9$���%��fΟn��j����~)�I%���%�1�D��(� �oeN�S�H����܈���I`�lT8�I���p�(� �%�1����bel�[�q �EJ �*"J��!��.S)��������Y,�/��X��o�+Ⱦ  �M��a����� �����bn/���O!��������r���	��K��"�7(C�}��1�2��%�A����DH�ہ��h���8��1=�gz�<�%�Pl�=�;�\�*9�K�
bP�!�[�@��-6{�/� �P�����O�a���� �-�?��|��\��o'7O�	�AR���! ^�h��H��$mcN�Sůs�p�� V�@ ~����y"�6uW�� H�J�l�$� ��3�D�X	�U�_q��	�a�0�=7�ݷ@�I�3��<~�I�aq �1��V�^�M)�O:@���/�y�5���� 	����3��?ok�sV�*�m8�Z ����(J_���? �jN�g��>��Ǯy��{�	��@�|�n�)ۡI���#.3@	��	zng�{`��D.(]J�� X?�9�Z-(����m�5C�g�:�K��Y;�K����>��%���`��ǳtIa�	�p���� F�v�������\�� *��������� ��0����
֢���ѹ�R���A��xV���rXIw�2,��5Q�������+���x!u����0���	����%���l����PR��N1��p�/�7�UV�|'@��\��[_���D�XL�8��P[%�OR�ᾛ�a���-/��V���8�%�����1�I� �?I�����v�N9���D��N
-���4e��U �ʾ�z���0[r/�/$:����j	���y�&Xw�P�e( H�hP[Ig c�����j"��.Mǥ�%��d��$�NL������] ������%2�� �i�a3趩�hW�t�-�������P��#Ҳ�]ؼ���a�ݰ#h܄sZR��f��Z�ؚ_��#�l�M��W���	f�v�y=�H�jUd'��E)%�ti�K�G����k�Z&�aP�~�Í=�W۠�q���t���%�8YqxE]�pH�Lk ����V�c�ׇW���\@��B ���g�	�s�Q_�]�'{�pw ]��
��Ől�ja���抠]�5��r��u.(��ν7L 7��a�����WV�I]	�o�#�2�_H[6�����~`����P��q/Ҹ\���}�HN���{�P��@�W�1�K1���*ژ��y�:'P�8sn1�#���K��?��z��uhIF������*�Mgd`-ڙ�|�M椾�i�[-0U�n)��:�揲05� ��f�+�U%�eX��@��U�[ {F ʺ�K~��.��Q���q,��z���(��{�	�Q,�!	�ax��x��at�1�A	J����N�N	�|y�K5�xA��"e��^z���)a{T��O�㰌w�{yJ�����^]�FnFER�^��eF(�<��r����^��+2�[I��8!<�Nn�~ ����03�yJ������J�� �	OW!ȟ�pA� ��N�Kr�j�!_��^n�>��3��@�DR,Q
P� ^41��(�p^q��7�����T"d��ҚV�!��	?�t����E))����Awi�:V ���	�
X�H	��YuVD`*��g'W~ESn^ u�I����%�̘l	��[\��59��	�-a��;z`��%0�:�K��4ךk���A�"�$$��o{!p|�����=@)��1^�C���� ��wC)�ؘ'�+ѐPu�U{[�<{�"dzoc�vHM\�Yf/S�`Y�}
5Q���__j��yo�
��m�21�=c	l	�{x8&',�BWu�W�R A=�}��I9/)�YЍ�`�Z�yK�͎6��XaZP �s�����o�0	�!�y�j���=W�5�%+�z%˘�uR)�i��]��m'Qi	�5y� /���՜�\�L���e�l]�`���&��JBD�P��)$��� (SR�ͭ�fN��N ��˚�H�֋g\p���*����q��bT@a��'C�F
���;_����0�� E�$-�t>�N�2�WPR#} )�! �_Z1#jP����^���_*W��:q9����nc# 3 ����	ɗ+��M/'Vf�T3�x)uz	��j��"� e��N��4���ǳ�AI�TB!!�߰d�.�p�-�U ����q'���L�:]>b��u��;��'�`X�A 2!��@Ma:0N�q�ɚ��E��D��"+ȀE�� I�ѻ��e��2	���V��\xG�H��N��[���H����J��KvJ�e��v*j4%۫�E@�������(�fdBA���_�[�A .�Z�;��Zq[��@(���T*$�H�!(-]��K�w�A)���6�B�W�<d`,�o�	���DO1��K[�w'+��cυ ���� `��?�p�)��a+[��b����e_	�̆"��`�=�`N9�3Y}�0鼕5
 �^�SI�)7m��oy� �'b)���R�ӄ]�[2F��@Jz� 6�r?\��������;	j��^L^�5� i�re���4`� ���@t^j� �i���˾Z ݙ�4��wENa�V[���%]�]\ZR���T�|����Δ�?�]�� ���W�]�g�8 Cx��+W[��`'+γ>G@�L�"�եK4�O�HJ5�/(3���h���JJ��1��k�jj���#W��}�|Y�0�ce�ZT���s��i��ɳ�/%��
����	�|1gd��c���ۖ)��;�`P��d��5�RaV�Y�E���U�ǰ�o�����m�9N�y�h)�'�Vp[���d%�#7H
�b�wh������`�"�(q�[�E#QX/2�P�,���ڴ�Ϗ�Q!����uo�EV���
j`�!�� ��u+��<�~���tI�  �j�ֳ�Ӯ��2� �N� ���"!�� $�D�Y�Ъ%	�q��D��f�[��V&"p�����i��_��ך�����/n� ��w��J)�e�/k#�7��t%Xg��@�2K� @����$�\#_���p@<o�J��� ��$,'ė����	9*8�f ����յ; `ʴ��?�hn[EQ��_/C�XZ�%:��ȷ��F�PX�wyĹ:�(�9O_�o�٭�����3�q�5Q'�ao)�ۀ!
u���.��ݗ����@���n����bM]����߀�-O� Z锚������	k�:�Ϸ�Ȍ�^�Q��_1����e�'��%��*�'��YȆ����]R�	�Y�Isepj��p+�wN,>��P��҂�EߒzQ� ���Om�����a�ĸ���C�I��-:'���J�{�l����Tبp];��ܲA�
�I�[f�ȶ]�'���y#���_�'�(#�� �d���1�}R��
��b�p&���O�ZSU_�>{�P�`��U�a�@�J�hF�p�wfF�:�|ԝq�����3"���tR /��n����W�5_:�K���)��a�Q�m%fU��i��x�\?Q`>{�;�@g�_i���e�<�g����9p`���,��11����/J�d��{�%���Y{K��v ��z���n=���:���-�G�-�%%�R���3Q#����+=+����݇�K?�ż ��B92���)��^�Z��/�\��&��pf&�������Y�@�Q�w�1Ĩ	J�H}�� �'P(c4+���4��n���Lg �-	j7���d� �%v Lpa��O]��H�K���sN��zڮ G3���V����aM�����cKq[� o���' �~\P�H<�|��� �?��e�X	�����z���@��AAS��k�<�ч%5t�)f�&�	Z�.��c�����a�[\bQI�_o�g,@w��-%���$�j��Pi�.��)�M/�@H�� tK�?R�_c^��	T��[:��R������h��_P`-����Z��K Ǆ� �}���,�%�%�}=��.����c�� i��W�T� 9���R�?G	n�ũ�kh��%_�T_o��I�S��KRN�p���0&ԑ��`> �������)����5�aq#/���<� p����h3`��i�7L��a�p��
�	�X�KޒC�"V[\B`�+. �ѵ'Ko�6(�� ��Ps�_4w��`!c�F�K��H0��p֕Z���e��	k$^�D	@�6��? `�F�ѿ���P鉸���_�!n �́ '��A������9�`b�I��K_�n؈�cیt����o%�?�gpM��Sƈ�*��j���ê�Agl��B6��g?;ʄ�S��<�M4�zG���'j7ׂ��-\s�5;�vm���%8��af�B>�ـԩװW����+��� '�}�p�������A%%��d)X1�-qӥ5�J6��..m�9{���3����%y��z%��ģ	���U���P}��������/��+�ւ�e&���\�%���ֿ���㌸]�|=̃�˹jF#1�<��I\9kS�p�i~)KS���J��1)���Z�K5�G5�O���A��K��Y1�K��.(X��v�o| }(&ܟ`��	pV#��y���[�z��yCm����>_)%�� `#�]]�;�B]_��\���%�h ��Kʍ jT�����%�j؛�-}s���� �7@;M9�� 2�(�U�-��o#�.���P�-�s+��#�xh�z
pٶ¶8t<�Tj�oK 3.Y�1�}��h�5F��>��.��d`���a��Z�JO�������"�\�`�R�D[%�	AU0��ߕ��1�q�&���Ř������Z��8���R)��A��O�]��I�`1`��<��3$��(�_C�-=F3�9���"�����B��%�ZR��o�Uy\��F �*g���02cF �.�0S3 �eCךh��f	m+X������c]�j�MեE��L��Ј]&'��w��^�`��Щ {�}F*�L N+�~�i�`⋟�e�訽Q�}�l� ����f�?�a�r� )&<�J��J�8OJ��m��)V�Q'Q���<~���񬧮V�u�~��z1������t�����@��K�%D|j� ݪ�,q�s����0�������`o(���j�/�ؕnp��Qy �4��������Mv(��1p���`�c 9\n$����r�_������1�	���}~U���
�� 4=���}R2�4eV^'�ϻÂ!X�:AU ��<����%s#{Y� L����
;מ�-�J��tKj�
�Q��:b���mB�)���-l/jbP���!�>�K褀�� AI7�X�M
	?�}G��u�e���[k�d����̗���i%:�ip��-�yHj�HC�y�I��/0#)�-Po�	��W�<�ә�?��+t̚6˼���9P��5����A��ݿO�ZU����&����ڢV��R�v�=��_�H���ɋj�c�y��j�c��K�C� .f������v�a[����J�o� ?_���
@�ݝ�%-.�l���M%//kG����6	iV1�W� �F�m!��E���CW�0��'W��<	Z�d��-ֆhT�i�.r�o\�XQ��_���ˋM�7� W'<ȭ}���.�`�D�}	X=��1�%a¹�O�`	���.���>� ���>>��p(#��K���� AC����f���_XJHH��"�ٜ �Vr�+ k�3`Rc&����" [jϐ@gX9��	ؤ�u{�^����ٸ����_ W�~µ�*��.P�`!Z����,��WP�DV\��7}�R����U���ai�^�*��M���}���~/��iT���OD�M��%T�Y*�aPJ��j1��~\���2�X->�X�����K��X����y+] �=��� ��b8���ŗ5���&�@������H������n�٘Pu��Z'�Wڈ�� щ�^�"�%��t璐�z�# ǳē'��!cŽ1z�%�=� V��)�� �m��b�|%)�W���t���'�A�7v핒��G�4�����y� %��/��0x�_���KW��uHE��Z�4��� �ov��m�p�Qڠ� � ��l�m�qK����+B�V�@�W�)	��6Xq���a���ûmt���Ka����%	�"���9��j@գ�.@ H��w�X���+���YxT��gJ'�~Ē��A�!�<S��4\����RJ�=�P��LZ[�ω����� ��>9���P������Xbzl|\��%>��%��i@ɺiT�L�t�ul=!����n/�v )@��7�����Z;�\A/��<0-�p�	�e/l �c��,n4od��׸I
/ Z�J�}�Z������M�,��8Ҁ��"+8��O�&��m&�L���xb� )��`y��6���#�^ ��	GH?Ҧ>�½y�Iaq} ��$���z�,��8[��u������M�\�aQ1��-.(Y^�,�"�2���/a�>^���ˍ�GE���0؃� �Y�bK�v���ct���n#E��ʩ�K��;�Ġbs ��J�[I�^"����u_�J���>� �jk6гcJP�# [1��N2�]�x��z�GɴS@�ya���.�`�m%�V��Xy�����2�)l�����"�)�i��kͭIy�*�[+��G+�a���EtYP�$E	j�tJ��$���u=�u���h���P\���?�ˀ�=s��h��-��f���0�9~�
�;�D���҈��OpT�1��F��Z[暲0�P}������Rܱ��w�Mu.�1�-is��m I;W��� �oi��\C�R���è��Fg�ǻ`�Vtz��m �nkqFXP���s_�U�삗�{#�{�i�[���<��^ہ(e�����U ��h����`*(�e�[�h �a��`3�)7��}�)�N���}�䈯"�c��"l �eY��[��3��U�lb��� ����a���%�`v���@"[N��V�_�6��n��90t���� ��" ��x��a/�F�T���ϗ�d��� ����%�
�P�[��X�� �[^�,�t ��mp'u%%F�m6C`�e ��F��>`L�'& n���{�*�X�$����"J_^=Q�P�1��K%� 4�&�i�*����&��u'�TZU �����1O��׋^0ip�J��&�20��/��iU��A�PS�;!_������u�|0H$��ಬ^R 'w�(�%+��`^� �j\q��_9O���E�{o�'�v�1���^B��?���7d��� ����ĊQ����;�IZ�5��k�����/ ��y��	�ӱ)�^5�윐�%����\�O��%���UM���C�[ɽ�J��)��������sp�)Z r%
�$K��R[����\G�F =zK�^%���_�C�t�'\�u�jn� �s���3�%�2�+J��%����.)�{�f��:\��RP�B���������+�g��%�J�.����V��^r�,Nd�~�?�p\�Q@���&-S�Y�~3��
�&�,�:�1���u ����8� �}N���T%�5#@�e�U(N$�I�o�Br�����#�D�e+�ےQ:��*�8vmO�\ZR� 쭹�1a �u�!�p}Vi�1��ZX����z��K��"Ŭ`-Pn�L�u-Q�b�ձx���i �a	DW�޹�Z�_�sQؑ��:����kAŷ? X�<����Kj�����	"� � x��m�zo��,�0]�SU�㞍�	�z��@Be�8����s�ѭ������+����_�{w��j��� PQ��J-�p\�i�ES�ǇA1&[/�9���'��G� %�[����%m]�[%��U�`��xia)�uoC���	�&�k�	�2\��	$�:�P�4��,	�v�����b�ly�g@%��Xo{	qQ�vs�'�T LE0�U�� ��m�c�M/��_j�2��N���L���A��j�v��iy 	qm��B`���j�k�-���z� �_����^	~��{�3Q���U�#Ɨ���H�^��p:�*"��+0u� �bv,���%����U����$k�-����+�]�t�g����4k¥��KE��Y	��^\���ʫ]��:�����fL`�p���^a�e�)����-�~Fa`Q_z�1D��B'�v�
��j1,�j���G^Q��[<�5�e�0a�5���?�^b���M���}U&
'K,�
�B��_� �>n} �2&��3��'Q��P)�S/ pTF�A��o@�[�	��_��!~FxE��mu~j���ړ�5���Q��.d��K���%vPYd�U拵E��{N`�U &��ER�S�� �c�� �Յ����K^���a��' �/j��GDf�3�5X�e�BHT:EAj�Iڗ�i��B\xH���e�'fd#��:�]�HV���Q39 ��B��._���U
!�MJ���D����a[��1 +�
��Ւ�ᖥ�hwX�=� ��=~�t3d���!�G�O>�~�  ̺�O�(�\�d�[�*̀l�(��
�d����J�H����o��n�i1%�I�3��ȱJZ�*�i�&W�oP���%�\�rCL��"�R��I������J�H�}ڜ�� =�Im[��n'�W\�U���O�������B�J��*�ja5�?���l�����R�^/.X[�~�.t�����4�9�������68�0��?؀=9g���('^	�xO���[p85ޖ`���p��fXZ7�aPZ��s�mp��O�iԱK�"�bh�u-0+��v2�o� 3,���;�HX�_��$w����+�nxX��%A�h�Ӛ�u΋"}���X0�8p;���U�F�%�J|��2�^Y@	��"�Smu+��4�����'ϗ���+@���Q[q3D�P�����z2V�/��/FV�P)� qNR�������I�E/P����ͯd`F0�������ܒ�NKę1���^�؁���b�"bB�Y���p-���	?8�Y���B�)*�&�p������l�k�x���E�мqV���1$���R��P��Pj��J��������J>͹j� ��N�Ь�Y�6TUd��9�_�A,Ne[5���4�_��y�PQ�R?6���wֽ��+Sm["�D��!��i����Z��:E^�}����_`�K���ךŻ��*(�O�yo`l���BvyKP�����j�ذ��+��)�" ��帶�;a
�M���$�D[�C����'��<J���l)��@��&w�1��$ ��O���.���������r��4�ړ���} �Q��+(2r�Ϫ`{����N�0A� )2���qZƷ��y\dz��p�������V��p�!�̈�_��(�p��!7�@�0rf�usP�E�1�z��*����p�C	\�d��0������\3$!�vPѝ+m5�Z;��C9�9�K�祱�Q:�G!z�� q~����F	Ya[j�7O�U�e1����� �'�g\�FJ�\�[����&2E�	�Q�4��,�M�Y� ���3��e=j��! ���P��Ϡy6��1r=#"f���%e����;���Q��p�ޑ`�Q�Y�z&'r-��WK.�����roV*���*�ʈ����|r�C@�s��G�8l5�0A�;KX[V�@��߀ :<��-��$�N4 @���b�n�	f�/�Y�	�ӵj��8��}1�k�I�k��؅Ϣ��9\;�4�������p1.�����qט��+aK���]�=�T�?��1'�y�A	��T��G�Ǔ胀�����0jB7^��Րb��^}���y+�3�:�t�I�|?�ԁ�r��)���h����b%U�!��߷ڬ�PK�VKKT�`@"O VN����Nݸ�DgB�����NR�  �P�:⍒ 5@I��E�6���"���9�ـ� �1 �`��gq2�b4 Q_a���B��1�	�!p���+a��P1mnn� >K�`�Xݰ��SL���pڿ�Q{���*�%��b����ɼE���`7�$+������	*�a����>�$�+��7
 ;��n��M+ҳ�Ё
�xŜ'�k'[�x�mn�ɕV0۫0����'�\[�Y�q^]d���+5��m���摠��s�	��9���;�������y��`	`���x �9k��g!�y(�8U�N��ŰJ˖q���G�� v'^W�Fԧ���������O c�+V ҷ>_��[k�R��&���z7��m��}��.(B��_Ǧ eqDF\%���`JT�%v��R`����:��h ����`[���ba
�V�� 42�P�ѷwH� q;+4�X#�4�c)�/�� =�1�~9
�-�&����Y%�5�7���@��+�%�UR6� �N`��.auƁR�Q�1�%{P	����/��'��h�t�I�Z� �KD1��p �̈��P|{Ѭ^�1� �EZbX~�aT�w�I����d�R�\��R.TU��.t��ӣ� �ߑ�1���j��&Q-`OI�| 貕�H͉����x�%5�X���+�̸H	�t�qՁ^��gs1 O��<�2�م��^K�F 1ʫZ�L�nD�zX�����H� �SG��@� m��b�_���P�� ��팏��y1���PRb��`(p�*,�``L��b~P[�|L� �{�;�k��-9,[̥y|� ��r�!4N%�V}@u�Z� �|�@'��n��$_�I�[y�H�G+x��6�UW��ط�mۏ8UӤ1��Z��e��=�S�Y� {ƿ�zl�� ����JH���ݭ�����G�	�~Va��pr�U����ӽS=��t$��9�2hh쇜�@E�M���ZN���@�,a�Z������d��A 60JV�� �9Z^����"�ҷ��ak�/�C�1L��l�1��ډ�iK�2E3���dD�f��Y���#�$h_��,
�a������q�[.`�]��.X���#�����Wl��r`a�YiKM?D��Ɩ�`�c�� d�L�4���[P�� 1+�ִ	�z�SЦ�A+�!���b�ŀ�(���	�%���c� ��k���M�dg����!0/$k&�p��ms� ��T�s�;ᭁ��L���ӆ��D��p�� 2����I��y�쵶m���]�����4�oķ��d���.햼!0����9 �Ձ�ʙ/�z	��"\P�YD`f����% S<z�H��0P��I�#XKa�s����	�'�N�B0��T�/6e~Zٷ�����(��'�Ԥj�`82�*	�ݭB���R`�[�����F8Q��k[v��ո���g"$M	�.{	Y��L���C����ۉX
��*T�	E\\�	�]��7Q`�.��%^a�l��q�V9���\�%^�������5>����u�����H������ ��M��ݐ�u':P^*o�o� B)�o�\R/'7��� q@�8������l��/d�Y	B�d� ����$�\$�� �c�{��Y	.l4��.@��%`,���}�[��.�������ID� R(Ռ�XH����J�T����#q�����I<�Ȓ�a��Z����)�&K�x%h����{� ����%�U'j�������h ��P��<�g�{%[�p�M���1���S�i@�kwh;�,0/�@p�0>}-f\
p��M�����?�F�FS`)��X��zZ��-_��[���ZeW�ϒS \�`��$�q����e6���Z� s����=���H��m?��mZ��[��1���q9L6��k�K�ɒ�S��� ��K��U,.�-�,��#�^?�-@����O(����(�p����1�%M$�?�����q��#��%�2�U 	~nV_%ď�O����LiۊC���8^0%���1�H�1���N�'���Ʈ_`�۵Ka�p�]�B.��,q% ��ͩ^��S��P&k4u�GJa��l��ǘ!lB�X��ݠ?����0;՚� �Z�[N��_	)��\r�hy��̹_��؊�7���(�B�K�r���h�Lu �d~F�+ �˸,M�D%�3W���*��&)`�K��<��'������� A:���x[������L.�=r��IǼ�CM���%Ć��c	8\�ԇ���(�ʩ�OE�^���8�H{��-@*���0�90�dn,�	�y@$�	�a�rU����
���	@%))s���S�*�=w���#`�<3X��`%����qZ)�>싒���Q�Tw���d���.�)�^o�	![Ȃ֕����_
�8@���Y�&fgy���Uմ/(aA/����E���P/}b�k%i���������MK��6�?��߲ˇ��n�o	�^w@)� R�-'J�5�d�����`����2e�R�K���)��`2Q��駗�vq4�j_K��x%6�W���_	pb��@���0A���;����"%���6`K��	z+d�B�7�/|���� �͉ji�y� y�F�<���A �5h�Dl]Z�B�V`a_�bG%s]jfw=�������ɯ~��ୈ�� �ox }zn��q��skYH*� �g&�f����-~S���+D/S�����1��\��F ��Nv�ߕV�I��)��b� �SXA���J&�!�[��Ƀ� +/����N����e"ȹ	z(W2�]D�'��BDX�N,H��n�Y�i<v* =��3�k��%۽��j�H]�� �%b���+~'|F%1�^:�hD耑� �2�гLۼ�N|=N���n�L�+o
S���� ���E�k	=��T�W�7@^[�X��1��cz����T%6j~r��zIao�O r��yl�#��D�%�2�ʬd�	���q�FYX��Sx���u*}�>��H�{\�Cg [����AG��Ҽ��|@%�|㗔�ĵ�+@��w�%��Y� r�>��8�)��j�F�b%V_���~/P�xq'VaZm�`翉�'����iK�݃+j- �
��J���@?���UH��f�Ǫ1��*�U�-���!��x��d !��YaPQ_]�S��A�!�@	��d{ç5b�����h!�mw�kl ��E�T��Fe����YҶ�V��p����[��Iq�+� {���z����r��>��\�{��<g�������V��?�OA���Y0�[�z[� ��@oj���x��%�gW?ǂ�:sЂ�UŇ�mB�yb�}��1^A$/�����%3�  �H��E�<I�S%�^�;ˢ	�"IG�����M>�N�5q |���d�WZ�5o"���4*���'֗��ZT���}�(�>���'�3|ˠ����^���L1��?��8/(�+2��-^�8�.Ը�
�u� �ːUL l��Oٻe�ʞ$	A@#�[/2�)a�*�/�����뜁ICˬ~��85��י��0�MZ�7<���O"�A�� 8.P��w_�V}Ԕ��ՙx�hʀ�&�� }1X�����	6,Aƽm��&���'a'.�V����[����� �}%M	��`�<@�����
�	�#��k��Z�Ǡ ��@J���p�	d"�t9���Z
%pJ�T7��	����a�l�=ݼ	�0,ܛAsZp��]V �S[����{�^�CЬe �P�b`!Ϸ��8� G S���(�s�	�`[����t�I�iq�h.����xT�{���p"�63�`W1X;��[f�%s���%R����1J.ľ��ҬN ����	�9^����@�Q�jJ��亥�0T[)�&��1�u�@ێtO���u*����}�T������ ��ל_ #��.���;�*������v�W��{*Y�%H��ݙ�� ��T3m���g��/o�����F��Y�;p��	V׷st�RsP�Q��!�.����~���&�g�=��<��N��l�Ť�a����@5�1*�M���j�������d���j���%�7�R9! 1��/�qgDU=������p`b�hTa�bq�t�d�D�~�s`T����%)ģ���uX^�;܌@��0� ����y� m���
&n(N[��W�� Е2_+��31"o�*~����m)���Bg�U�t�C�'�g��c�	K:U�!�A"*�o!�"��NL��Bs���`�º�TN[� ��@�:)p/b���d,��b9ה��x�zX�,V���n��nV���t������jÍ���dm"�2�?�jY^��c�ͶWi�E�-�?�+�o�'��
����$W�J��i���s�-/}\dԆ\����N�$��9�p�(�ԉi1O��BN��.A)5& )��J�n�x�P��J�,�w��= y���h�m����ڸ��~ }����
@�Lt�~���y] [��:���@�_�Ҽ�Km��z���/8�u�+�v�퉊 ����k:�߉�1y�DLQ�IJA����`���h>^�'��� [k������ ��J��*���`�	��aQ�/P.�%�k >�V?PhZ	g�]�z�'[3���>][6��̛`�P��@a�����%��X�\���Y�'^����}�G���j8੤R?|���Hc�]�Qd:3GR[�W�<9,��V�ֳ��W�ajQ%$o���u!��`OM@aN��$q�J�%v�ir� |�T`��-�H�N �<�p.�O�%��.U��B�]Lt��f���7ݑ��@��&�Y��)�M@뿆�!��L\t��\(O�t1��Vn�E�9�e��L��^E�MT@��FZU�#��� 4rb�h ָx+TF�M^��ֽq	`������9_qv�ʦ\m�<���Q4|R�O�R��7ʰ�s���%	)�w�~�L`	��  ��S�foߵ/=X�a����JZ�/� ��6wL��^��o�8����'ѐ�ﳰwU�0���D	�V���`_6�H/'a7�?��iV���.��B\i]J�X�E
���<}���C\�[���_(�DDRP��{����$��	p�%�	"]�&�tC�[����� P��M��X���������"���Iq�D+@��;��v	㾜�<�43�]D�OU4����j1��:�D�1��+�Y�^����Fs��`��E�3��#�pWf�}[���\�Q�4=�b��B1�W;�{R_e�a�����K��r�e��T��Ū�.�ߩ:`��pc}�GH��� �yi5������l�'�Y�$Y<�����T� ')�	&v��E%����,����)��K/�-K���N���!^��~`s�GQĀ�	S0[`a��%�P�� �J�ֿI�4^�VU�:�n��%o��v~`7�pE�� ���BK6�j#�Y��0-ZSbءE�BJԴ`�a���u�h�i�g���������jawO�`�:nZ�ߣ��D[��5�_]��?@sv�#�䲳r^S`����RK`��ê����Z�-)}\�������ƅ�e�ܞy �z퉕I�����@����'Z��-	�aW�}^d��U�y�b��c�fG�[[P]�$�����3�� �.n��	3�p��Х��.�ov&V%�D�鉮�, �$���ȋ��g't.�@>rt���[R�����q��\%D�RW�7}d��������  �~��S�. ��I�y��NĨ����[����.4��ݥfПd��GuEu[Lz}R'��%y"��S�{IH��}yv�@nXRK �\~�p �����i[�x7��$E���݅�(e�G"	6�oc	I�'�3 ����Z��E
�m��glڂ~��m6LǮ�u��!/-o�8��P>"%s�Y�/����	��T����	'.e�e�P!�	�~��{-XU �Ka���s�!H���V��_'j�M�u8����	.��?q�S��p��:�s*���G ���EI��晻%����u7a8�H�HI%�8D'���ղq�ҁ]s��p��7��L[�I����Y�Q�~� ����]���.��Xb:�	p!x	<)��& L��8{��wr32��O�Ȋ9B ���v2}Uq%�º]X��q:��	��y���r��Qn�!hx��'a	�Y�h�qR���."�& `��W'S�"�Ya\��v���P�b�%ë����zO9����tB�����/縡�=0�a�1�&no�Z�i��F��ޮUN��0)�1��AX��a�5��Q��m�Zې0Z�ՠ�_p��t��T�%���.�q��4�O�	��M��W0�U ���o\Dxzd�	ā����]?����G>�`U%�� ͷ�A|�F��1����HaK_�1�� 8^��W	+��WNV�M@O{:Ne��E �U�0h +k�fG��D
 �XE4e��7 b�P6��H�l�Q����B]_�tvھ�z�3Mw� `·��"�K@�&��&�ϭ@����	�}��DtS�Ep��c�	��� �5	�% m���t�`�ۻO IaR��h�XzM�K�;4h0��KP:�� cx=�4aCs�S�0tQz�o(`�+?	��<��,Fe`��9��V�k�5��y�z��j����`Э�-9)��	�`�	����,ȫ� %��	�x���xu�H`va+�$s�ᗻ���[H����z���"���L5��?&������a����uX���< ��{��x��������܎�_F����!=|���9��~Q�!�_Y�����Kj����Ug����h�������Ϊ��S�P�mb�����=;($���Z�[�'�,&��Tb��`o� _��9��k'?�B��f��� 	6���󢥸ʝ���Z ���'CB�oGn`�^�N��`�1j���Ƞv���b�<��a��S���@ ���0A�	�J�\�1d9#��ө#�� 4ȵ��f�&�&"�x����ل>T�@X��|�Rf��lw@ǁ�����n���tZ��D�h�vB�z] �G����U�8�Q������$�ݑ��� �c�( �vs��>L�� �#,����p0ОJ��h<�b��{�sH�'9�V!�^���'-�s�=,�X�lh;��3��	+������桵d��s��i�1�	�*P�MK$��>Pp��:y�o�1��k!_�UT��F'K^�Q$
O��,�;Y-��%���ы��Sݿ��b4��q���{MR���썒-�eVd.�������2[����	q�\�X��ح�	D^��F-�W';^ejł�=�<ď�{\��٦�M"�#�P�)Ka[�w����tR`���<'rB.Ok��.�'��:��}Q�:$���eJ�	�� ?���h_�k*#���Ɖh!�MB��M@i��a�����-4J	��{�1y�s*12P`{�3%�Oh#_�W`U?��ò��ݩs.x;��ޛ�"VP���j[�Nw�;�q�N����)1M�4pQ���&3��qm�P�)<�� ���R
ء�fJ��$ ��n��Y��徣-B1N�+n�?��RX�2������t��
��Ǔ��b�&�:�b/��t���m#��@T�X�&���)�� �����N��7e�^�V�5&�	dA�Mڹ��:��>6t��qe��A�f�`��{=�����xa3�y��A����]S�I�L`����+�L�)�����2�Ȅ��3������I�b	׷��x7w%}
�=�s;'���e��e��ؓ�ν��P�T[�`(��@ �A8���Tu; ajד@��P[�� �׳��.�Ѧ޿	�Ц`'R�-AX�ABa�:(��U༤fY���`	���j�m$��O��lϐPT�K�|��*��0�:��m�[ ���!;<{�_����.r�p�GIlJ�R���+�nV�VZ�k�$�����sebo[�����J������a0x�s�t�90���� AY��)���z�{QK���	�*��9��:d6�ґ>�Ľ7����	�u:78������E$�/L� e�4����d����	 �a\�[V�@ƻHS r7�e�P<�G���E�^��7@��?KA;��"� p����q��m��0E���'�bW�q�Y'>����`#��I?	�%R�awDTK�г���		�Y�F� �dO�,�ѻ�|_&�X#�&��`:?ԕws��\�{DL�_�K��+_��	��-y׋������>|��[�� �	��"��b�� �\�K3��X�y�Ld_^�`����lmE8{q�$+��'��
�t~��!�` �\��m+O���at�-�Uy[��=/2��(`и���z�a�H{��V@�)�	��� a��O/�?��X�Z�v���ט'� [�B�H4>��8` /+��(�������������%'��MaI�.4ڌx� ���	��u�ޖ��>�\5�;o)��N�[3��~��L���A��+�	���l{a �r>�ͅp��}Q,���X-T!j]a�k��>j� �1��W����_ᰀ�_�ʈ�k�a�أ����⷏��t!㎍s&n�0�����~Z�� �%�CZ`n{/S�$��`�����%W$ �r~���$jP���I2��ը�K��M`yA&;��s>����~�"� �����"/����[���+폄��D*){��LZ����&_��"ڋݩ��LG�X��r��@&�Z�1��$���@���a�?�� I�T�N���Z���^��2E�.(����B�&@����	`h��5`�����	!���%y� �O��\=}�lx���M\i��*�A������>$$��#�1�uMTI�~i%4$����F�.�� �����1�=5A>!���+����h��~��-�>�ނ|	�ma��د��ܹ�����	�.Uq���1�Y��*W�H��v���;�}�L��ߑ@,ay)��%��t��F0gx.�J�aC�8�D�Z����_��S�'q���7;�Q3X�`0N����t=�Sγ.�8w�OV�`�̀� �2J��Nگ<	[���j���li `�Q{���^�½V1kޟ%B�0�Qj�̔0ZA��}S@Qf��|g�3H�Y��ż��<z�I ��ެ
�tg�	E����@J	�=�J���b�V\"��B�Pw��/��VN�8x���c�q�����C��P>��0�q�"_���k�# ���Jx:DN��Q���XWZ�E%�b�����s�'�I+���׺��B}�q�uE )�9�%�80���	�\H�M^�����@�*} �1�ȁ�TJ��$$Wóm��_+k�# �}�)	K�EzwǠ�����t�����J���%w=�q�_�0��c��P�� ,7�q� w:�x#�c- PR��K1��^��N�nP9� Pl�	.א/e\�޼*�a/+��j�>V�����gwJ���`3ݸ���MK�Ͻ�%�x�Pwu |��ˇs/-��-�z�F�kH���/��Tg��J\��L�Q	�,�NH��֮��0�2 W������:�?K�zRJ���m:g���ϫ���[� ��
�1!�\��2�|��Us���=K2�K&i3����/��"��q=�k�4�./��������)'�5���"�	l"�'6�tm�����V`���8���}Ƹ�:rF���|)�r��V�V�@N�yg{	>��Q���#NBf��R�����0��AB��[wp� �q�˵sh��AR����A)��+-�P�k؆K���H�"%u��Io�S���2������r$,g%~�ޝ\�B��@}�_�QU��)k��%���PY�U��Ţ7�����n�ƃ�����%IBl���� ڷ6
��%��!-��^;�L0����s��j�^6ܿS��ձH�ݵŅ�)*`J orې���0�M@�KG���5a�X3�c�	
��q	J�a�+K���Y�#�Ȁ��C+Jb���w���e	+�$˨��./���+�&�+ȉ�y2e�)�Y��"��d�;d���
��'�� �UCǀ�M���>PL=G��:��'��V*�E)��"�Y�NE> �k��q�=�рW�
��� �2J[ج�#�%Tր%��tP���k2���V��u�7o�R��̒�~���R��Y{��V%��ֈ�y0�V��{`1�	��j��.�s������@�J��u�����8�t$=���/ԝ׺�cUY-+��:�"�s�����3�$V��m�`>���-ܕPD�v��-��a#�Y�Īk�`f�x?ank�# ���(5�&�������q}.>���>���h���u��ν
������gw��;/��mv1���?���-MypĀ��%�j������̣�Tf��4*^E��\_Գ����Q��@�K-�,�,N���s�RMj���B.(�M��(Nʍ'+ �u�V���;�p��MxgH_����@<l�`�7] Ԏߚ\�P_������+H�(�f���Vǝn��,<��U =��� 9ɶ�oJK�Y�Lj?���{�-��#�G��wP̺� �y΂����Q:�K�_P&�"��1�U��%@h
g�֧�`��� l��#BZI���;�֘PHX�a�� ��9���q����@2[cyJ$ն�	�s����+�DY��l�����@C
���@=NH�~�"����82���\�a)�ex�J����%�G��]&`�1�I�X�% �
9*�+�c#�6Ka���彸�������r�א%�� H�|W߭�O��.� �O �5˶���$��y �wf�O�-�y֭dR�_�lx���C��/D�W�*<�eP��-��&Z@U���|O��$p��� D9� �m.sY���#�^�b7|����R`3X1A�n@�V���&`�����*�	;��j_ 2��V1�ŵ&ܐ�)��'T@��sD�rl�w��f�����%�I͘O�� �ĉy���s8`l{����aͫ���I��8�Y����e�X�(�cq. �N� קΠ �V+���H.9%���_��@w�˕%J֨�8�[��Wrѽ�  ~뉽�Z-�0�k' �N��e Q��1�_��*� 4��j��\����91��xN�.:�^z� 4~��H�6��NR�n���QW7���S��տ滰�J9�p������&����r+ܒ�MN_	�ɜ)/n�	~m��f���A��q!$�
���:����X\֎؝^��,'�J���d����oJG�_� 2���t�F	Ai�	�v'}Bw7r%��*�1��xƛ�/�JY� ��>M~�DZw˭.�����t>h@���c@7j'��6LC`f�Xޮ�,�9u` .a_N��؄�tx�t(����d̷�{�� kd*nJ��]�Y� /c�N?� $���7d9N_�3"C���P�߂�0�U�.n) �d���fmB4����<��k��������lf�!�U�<�#�(P����da�j��.)�+�ʻ�,��Ǹ��	��L7]:SW�������.	��{�����-Ս{2 ����J�	5�x���E��g�ϋ��0m�TL=]�F��  �P`���a�#���,g���W������iW���/p�==���:	��>�,��x� <ðU�`�	PR�dn�1����Zg��4��N� ]�4|.l�G"����� EJ�X܀�ӫ ��OC]j��T �Z!fRy� 2:�\`���V.5� o����d�l��Z�aU�־_��*#����H�!%���s��h(�AjO��k��;:�Ej��`�U�a�[��s���cw����/����G���j��?`+�+�f2��^�X:���/�b	��W�� ��X)P�yء�n���φ�Ӊ���z#{��cj�6��{������.�+�[#�=Ĉ�,%�]�< �2�q		�W���;Z�߿^��"n��"ם��W١(�����+i�FpM1� /��"�阩I�`iIpN$DR��7;[/=`� 9�R�fE~)�na,	1	���U���[�s���{U��@	�r�y>��qL���A%4\7�/�� ��9`�� $ǫ������T`JA�B�E�.aP.���tj�g�	Z ���l�_�{tr�o�Pn���%O���륛.�y� �+��p�'/3^SI�mt��IB��9	�/l�x�J.���e�ޒޟަ/\vԖ���+'��j�ٕ^hǝhr��P�1�r�[�B}q�q���]0���s(�H���1�u�/�ە�*R`	�奁�ܡpa\z鵻�l��/)��A@S+�E��y8hr?X��{nW⮍�G.��n�ڢ]l�xr���8.(iw�2�o� �<"y눛�Gj��k~ �0���4��`�Y2������.M���&��p~�v�@.՟ "�G��Y�<�4���Փ�_���4�I���j��3��K��� �t�	7P��
����}�Yj:��������h�0\H*��n3C�6n�ܼ\��^�e�k�5��S4E,鴿&�x%���3��b+aN*�4mۮpr��.K��*����~e�vPQ�Y�T t� ��i������)�P��{"x��VM�]�	�s��F%����*O[�@y"%3d��� ��q�i�^pa��+ϫ"6�� �K�M:��دD�[E'p�b���f\����Bg LfקS�$n��f�i�[X���KUf��߃���{' �� |f"�.��f�woY�@�&�Ln���[9^��P�������UpŽ)�a�	޾Y}��o@��� a�5^��J�#8.O���;��l���!#��=�J!�=����Kk�-׷p�ns��*�p	�{�`J��"!h���Qss� ��u����Z��q��"�'u�1y0�V��9��s��1gub@	��,W7Y���%�s�<�����q�+�d�������P��0°c1�nH�7��|���j���8�̺�t��%�M�F9�1����px��g�{�Y�'1�\��p>%%n*��%iַZ_��`V6�&�p-�!�d����q)��%�Ғ��80q'J����YP*���qC��$�C�y� ��v�"���U��?!�W<���R�_ف���V>9�$�Ͻ�w�_��;:�"����1A��9.�9��n�_�v2a�yv��,�U7}�t���'��^	�q�jG����s�i ���O��t��y��_j��Z�g�� �Q�B�ulE��6 ��{�%�r[z;E�=$���v �ћ!w_?�sڱ���������b��U�b{pa������g�o� ��������%-�XB���Ĩ^�� =���z�j/�<TDj�eZ��$ƞ �MP����'���l�����Frl7[:6Vy�!K������<�or�I��@��%)�}����ؼ�Io��`d����lp�Qa��H	�m|�I)�>��J�h�0�>��y$-\�8�P����������+-F#�=0Ϛ��E@�\��z����)�a*y��ڔ�;�>�/��~2�S9AZ �T�_��џ��'z��%�g�V^��QjZ�{� �R��4���g���?�H�	VQfõ��ۻ��O?S�K��̢�	���\\Nqz!�*o(&:b~��l�����Z�x�E����X'�tտ����'����P`̕���y-���&+
��}a]}}X��m��`e��H�F����*ۖ���\�%չ�)����u,��퀹�}icu�%s�1	�qD1a	. ���1��+���U�E��1�{M&j�8	����~�-W��+�`�f�/1T�Fan�|�ѷQ�E-��oL�����* 6Ri�|�<��O��	�qZ�&Kĩ�"�~�a��f��[�M�qJ{`Qɞ�K��E��#%ג���'�0��M��lr*�O���9��L�^�T(N�FS���U�����Ƨ��f���B�jO�@��	���7�[JY6 {3�|��[��D�z�v��k=?U�!��u�Q�`��y�`�!�	���p'W ŀ9d˘�2��=)YC���<�%��'H���@YGj�����{�^�@��7�='d�xSb�Q��VjK�=&߱3��+�Қ���ȫ����]#����q]FdD�͡�L^�'�/��u=*
!N�����.4a���!",*���>�VK��O�������\<Qt��=j����f�%jt�V���p�1q,ԫ��`�0xg5���F�����pi��I�x+�Q�[K�����.���8	.KaD�Q��O���f�d��!��~�%Fw��>�tK�j� �^�\�1��t�P��0pF[��=������uX4N�(��N5���%[1W��X�Js�5���BP��V���B
�~X���s1Z�y�g����J��{$��A�t�n���0����7��o�kr� ���q���=s:�Vpg�������P�>�t��J��T��E�`7Ť�K����J/�����o
# &5�#?�\��&I%/�#eF���)�q�����S�n��a��x�YŖ:�i������I	uμ��x3:�h���A'8�tL.�v12M�% �b=�&�$�,*�� xQA�p~�
vYZ@]�%j<� /�&ё�u.����'ӎ�1 z�wL�����c��P�2���3$���W��`P�!Q�u9�S����Ua�<`��X���a�UI^ts�N:���+��$N�d"���:�(NF�_��N%�;W����.o3`8jQ� �O��.���ڣGrmm�=X�-�Y�%�L�pcF�b���W��]�� 
��_�Y)�G�@.W.(MP�s�(G%���-���E�<v9_A����z�����_j�)�N�����&�:FR�=K�(/	^�8Ć�n
���_[b��wؘ (X|�nB������*�|���y�욓������2Ih� ؊�;��+���X�K�8_(P�VM� X��J3	�%^#�*��I|m0�eYP�/���c3��#�� ��v�{)��%�4��3@� ���/��UhX1�i	���}�%�^�Z� �'Z/�_"�9���`����a�f	���(}�ݒq�)���ߘ(}���Ay�)��? *?b��:����s�3�Up啋�Uo�d�ĮZ�j�^`:4�ȟ�ֵt�a���8$%[�S<�������������4S���%_uٻkG#E��U>1�.i�{�j{
��)��������3%�t�UQ�5.�u_� b7 �an�кZ*�i��/)�:�t�{�`ܱYz�J�xJ��Ë�֍@�s���+v�t�_�w=��С� 5�N"�����������ш��v��,�x#�'90\��f�5LP=���Z��H����Ł��EM5DX���0	��W)�����/��oPVp�T�CK$�}j��x����|���h+� �"�l�w�Z���������K�@4!��zZ�р�Ȫ����!c�b	{O	J^��j���(�P��2�K�!��.�����t�ԄNX)�#|m-�\֟�����V ���/���	Y��3׾��� �|�5�����ʰ �]	�$�R���ὤ<���r:� *�G�d��v�ͨ(����\��W�Q f�G�a�%T[[̄�)9;���@G��[�Л���ǈ�0��Oc��/5��@���1�:	���Z	���'pW�3e[��r�	�e]� ���݈�r�dm���H��!�ߺ�� ����r4�&l������� �^�!������o�t+���3��ҹԁj^�\�R��_����ᕀ�UGI1�ֶ�`��VY{�*'	��Bu[o	)�z�(�o7}�K���u#��(\F�NRȪ� y�<ί�+[ ���*�X�(�{�K_� 0�=A�$�����D�K݀H~�!���_���	�}��p`$���mI�a�m�D��� ��{�]�	�2��ݢṶ\�-��'�~`���rLo�,��[f�pm�"�^�����kP*V���ϓp�c�X�vpB+�V�� `{"o7�-�Wu�˿6*s[r�N�x��X��$~G�%|Voa�-.<=��l����'/qB.�Q��O��격�9&�7��b�WL_��'���ݫ�J���_�y#��������	C����;��]i�� {ڧ|�תn+��x��	��y/G_i�\� d;�0Vy��.DJ`�Y|�f��qa/(����#z�L ne'`�V� 	q.q�/]�� `g�0 �k��_Y��a��"F�tHM!>����Pҕ���!�\=^�骋���/��yc"
 ͔H�^�!����[�`k�� ���R���3�ۻ�'�S�Jˡ���h	��e\dV�{�Xp�)\��O�(ڌ�;x}^�ȭ� .8����� �~���v�5� �[���%7�<���_pb�	��%[�%t��!ո�c�%��*{���v���9R�����V��	���-��
��!�-��M-}�\�ֳ����Cٗ;�R�Z-9 �6����$EP*`�#�6 T�C�<�p���W��`���Sa�F��	���=qԥՐ�D�	r��n�\�z�KQ����['l,����Kх��,�.j�x9X��oy��/!Cw�	�L5�U0�q�SyRM��3���N[�H-%\:e֮!�@�}2�KKX6���7�#y���b���7�:YaeMb��x*�LL�şW��{B#%qd	A���T��t�	��vS��6��]Z���D�`�!�YT�b���ހ�8��	��n���yT-w���y� W���@#�'�Vvq���b�)]��ƥ(�t�� ���T�Z1?�4j�1���/�	���\�W 6׷�b� �������ZM��;��%�ePR��Кz-v�S����%�Ƨ�ZU�0�7��`�Xj�����Yv� ��~���P=I��� A��G�Ǒ%?e²56�(}l�X� �d�#�v>��}q�kM�@'�AO�"�WM�c7��b���N����	�W��X������n��K��{�tЦs�̫��ܫ��U����
��Y�\ 5��\!rM��a�W��u��EJ|� ����BxOF���ě�q�-M-�OFT{ƌ�1������� 3C�]y|�*���>��a��{��x��4�@M`��̧nx}
<�UKu����߽�MF��f��<���JB-�ٿ��z@���s�*��է��U�z���L^7���$3�mJ%�� ���^k�Dw������5���!�v��������p�	���g�b`ro�I��.�m -�>� T��|p�k,H6|T�j?���~ �)�Q���r^Y�q1� ���Tu����Ch ~��[�4/���X���*�����H�+w�W�P�������41a2X�Pf� �_�Fxn��h��v@�*�� dv�UZB���i���{��׈�K����0�� �E,r� Gyf����;��C��-�'�X��G�d�,�^�)�ȝ��x@�p9�@��=u��Q5s "�M9��C�<!���^�Z�� JL<+�N����{D�!��Ʌ^t.��"�<7��X�ȸF�����1 �h�F������H!���07k9�^ή`Ĩ��4p�����&O�\ �BW:1��z�ܱÙ��s �9x ��Z�~�%��X'�!E��:� ȅ���br����4���jղP�;�������Ȁ���Sy���F�7��&�s�!�߸�O \pF_x�m� �r8�Ѕ3Z��(覄�ɔ�@N�$�dlʕ��Í<�!�d��;�րa�*��Q`M)�v��P@ąp���B�~C�9�  ��^��%G*P������N^ P� b#�J�wI���ƬW�
}C�<K�^�H<)����T�Z�q��� ��ӻ�	=�+�� ��� s�aU[D�1 ���p׏3
r����}|��J� �/D#g�V�\�ьs(�{* �	��ٞ�� 􄹂=�̻}�;�?��L@"Y ����1�o>t[��G�����A�ؘ	M!g� ��>;&I5�n���B�[�E�	 G������&�{�>���!}������YU� |����Qa[0���ɰ��?S :K�[2f{�! �i����#�x�=`_�r��n8x��!���.��� >Mȟ����)B��
�<�0&������&F�"� ��P	�Sf ��>a��P�R��`$��}/�{ 9D�(���v 5��hR�� t�y�� B/��>���
��H�`�@t� k7>z��ۡ 2��U��\�)�V�<S���Q���������(X�o��W���0� [���e3��� ��\�`uۉ_|9��vH�TB}t;cgmJ{�dSnUN y�=���'ؓ����`��� >}K.|-�6W%�c��� M�pC}��6 jQw�d�$(c�����;�� Mǹ�|i� �,��c�� �8ܟ�D<p �=���F\� �+��a҈ �,�ώ$J� �Y<�1*p�&�8��h��_���' �^�ĴPSX�v��Ȟ�@9t�8�����������Vy� ��X�m� �#�s�Î ��"���� ��!�ҋk��� ��㞍@w� ��6р�>�v�L���{?/� �����0�(�-��� 1���(��{ �U}��T~�x	�k
��.d� �A�����,>����I����L��l�� ��3����<�V�?[�j��4�p�8 �e	xc�#{`!��.�~ ��<���G�5�E�����F���˞����5�  _JS��H����V�4ԓ&<���C���8���  r����� ���E=�j�ަ ���	��Q`^�>S���ۘ#D �si@ho ,�Y��Nl�H�0	n� �bzQt )�ќ���w �|�?IXJ}���n���%� ������< U�=T���8�	E���� ߈���* J�>	����?\��Z}�sB�I� M�ֿ� ����KR� 0	��ɧ5@�BM��*���	 C��ji���5�$ce�s��#'Oha|HX�;� �tS98k �������>{� �����z�;����!`9��y�`$1��n=��&qt���y��V?<.r ,��Q����YtzI� |A�8�E>C(�y����td ۥ��+D�4 6���g]�u� ݱ������TF�t��#  p�l��Td$�';��}�*� 4D���Ʋ`i~����w$�?�����Z��4���C�A�0��E�0=6&�c�`� -OJ��9	�R  9�0�{ ���;'yuY>N�p@� ѷ�ǓU'�,nI Aqt%:x v���j��� L����4�iVd*���� $�"`{� �ѐ
�>;��� izXo�1� P9�<V5�=We��t ��S�y9%[ ޡE�����G�zq|�����<t�v��(��*a� ���;~��.�RH 8�ȪV�Z!FX�(B�<p�E��w�x~syGl��c%��y��5!�������4q!*\" #~Q�!�����s$��d��:�I�rw� ��4E<��p1��a���YX~U�8������Q�f1�P:F��yz�4��0����}xD�����)&��@��v��
��� �E�� �\1G��{�9y�xWy���U�$%d��x���~���N
����"�O��H&w��e�,��|_�E�D��4�<��I?~�r�nQԐ�P�X= �l��y���&�@:�� AY�@D�i�.�3�����3 z�M�R%� �H��t~�b㰠�X��i/�X'�$�`��|�f`�����~����X���Q���� &Y�z'�o|� ��}�� 0���f8�0n�!� dl�wy�~�r�䛋K�x�s�J
MgR�^g Z&Kn�c�a�A��ൂ���_8�!~�ӵ��R�y��qL�W�/�	�*G����ec΍�z �nj��y
 �L��{�|��8O�gލ�xA��;ˀ� :	R����p��t�q藝�~�'B�|��o� Ӧj��	w�6�!���c�q� h�6��b��L �~�9���Iq���R;@at�H����p��;BO��}�I-��"�W�v
�0��0� }L<|0D��X�V�135 ��ڰ��j̨!� =/��
�1!ȸSy��0v�pXJo Zc[�>� ���\���Pۆ�p�Qz"���.� �(��}�I� 5�F��M��@��z� �Q\G, Z��Rd� [8�_�n|=�}�s^0�?x�,�-� ��ц�_�c�m�f�,ǰ]"X �56.?#��֤Up�4 &�\(��z�x7 �뚔M&�1�A0�� >��y}� s�;p�ƛF ��6HT�� ����%�9 �qN�5ǯx�~~��r>sgk��� n1&WOE� �$Rs]%0����
� �u�g�e8��ռ0�( 1.~M�6,��ܥqz  D��v������n	w��C��A�.t�ۣ5�n\�� ��O�e0��Ag؉���Dz|�o@IA�TKC�o�ш?i��Cg�P <� ]���v�z(h���W)OJ_�-uw�Cm'̈�!� T(�/^� q�ri�(�������� ��!,n��+x���?u@�`�<y ��̪RpT==r E��K�� ����H&���� �s�u�t� /WEP�� ;�%=��d� ���M� &eLꕗQ=�x .EI��=/(��Z��xc��7�T��|	y���}bC� bT�$�P���?d�c�0 �H��ՀJ�qu�0Gw!���vI�P�M�'�9%���������(�p1>hx"? �b��T��.��y1�]��g�`�Q�"b�|���� ��:���E���@�J Z�����bP�*'���Ր�� 0Jӿ-�?�t���Vܳ��y�TwǠ��z d� n�k�` <��1����r�柈#ժ^R-J��9��M�	�C�� _ �Q8d�С�̜��0�N�2:Dt'���������� *CL1 �
g�N�3 �#1fXϨ J&��<�� 5�����l ]�\$e�U6� �y�E3 �%*���z)>��:����4{��d#k��H0���# �ņ=��6��R�?����ڐYg��U;� 홰�	s�^����d 4��CH7��u�����:�=vj FAI'|QH��!?Nim���x"Eb �!z�y'�  r�#{�� �BQ�"z�c�����p(�!ǋ\��m��|�@�sA�.3�� 6�xݎ& ߗj�+W��o�#H	[�0�� 6|��j��]?��Bl^9�f� �� �H�� �dL�=%�	���� ���' �,L�i[��w���~W-^ �ʦph�/ n�q��CE� �:�Dd� �%�S� �U��V��~,�*|e�!��s� p�[��h��ե|�P��Xƀ���Dc� "�Pk?� ��x혔�A.(��0���Z _�K�@���x8d��`)��T�@q���0d����*�]�H� >�������>���ˀ����=���f��xC��a�Q�����F��:�2`E����SQ`�I�F� BM��gw����� k�P�{�<��u���k *�2�Y֒�&8I� t7�~ R��_����;*�y�<�� 4ƞ�8?�pxE5}0v� - ������bu+,&".��gq��OLV��^�r b�gʴ�>�M���r� ]J����"� t�~��[Fl�6���fܺ	 �C�cs��Y�F0-��v�� ���w��X��B��o�yHqZp� XːO��S���`
m5�R�Nɵt�?�C�k� ���zu�<W�y�L��P!h��� �B�<�� �Hg@���� ��[�j��6�(Ƃ��Y��؛`���kf�@�>C?h��7�������fy �%�A���q ~ֺ����]�[�	��  vb�_�#� �s��lr�0��(6�j3Kv��=#`�!�B)\ �U�}���@S˾�=�Wv�8�@�L�0� �{��`�a�h�(ϴPF��<K>@�P���A �,�'��V}�`�p�S�D��;�/te|��k@�� *�9R�Ck6x�t���G܍  {��Q�?��V7�LY| � �2��i �b&�MD�H J���S)6p���P�e|`=Յ�*r��7����?3�
b��Ʋ) !� �`)P��~ ��R׏zx��\��<�����A8=�]�S�@ Jو��4�}��f ���n91�!�������� UJ5ojr�� hp�	Q9�O#x�N(��[ ��q�"7�jE����*���b �y�֫��>���&vp�@�h�LK|؝��1|%}� V��m��� ���(���f0THʻ� K\�GO� �AX�5�����#&q�H���f �4���� 0��n̓Z �Ag�W��� M{z
� E�Զ��!5 ���#�A���� U H����+N �BE��<�� F���t�^�PM�G ���P�� ��uO˟a �;c� ���H�x9."�@;߁`t�> 0\��S7���E� =�J ᮥ�s�M3Z׈ �T�%� z��Ұ��f�X��@��&V{M�UI ��u� D���հS���IX����Z {5��Kr�0�|���� ��P�e(, Zi�B�r� �W����L� ��E��]�#���C��~�`�� �g`�x� y�Mڇu� ���ۛ=J���_�)h�@$���$˺T D�pƄ�]"(R�- 	��y �+?I��i�0d��H�{n�� `��Z��s�������������`n�yFi�҈%aoB�������f��`�%@�X�p 8I1 �/�O� �)�?���x�t���:a��m��� 3�ɖD�nR��t�P��N �v�� ���}.��: �#�r��h
�� ����v=	ŊT�X&{ �\δ?�w�[�� �l��j�
�t�d��8T֒�� ���Z�j��3�p������ cG����3C }�D�� ߲�V�;�� ι/޽�I3$<ꩄ�䀎A�R��O'肨8��T�/`�HS�$�ȹd� 	e�o��O��鏀0�s k�8gLYnm<��� ��6A�)���`�C���`1>�=}��X�����K fF���E��y0�����+Z�L��Ρ� ���b�� �w\E* �1r$����5lB�bg ��HF�$�҃���- ��EM`�f U(�˫�O�c� ���������bbu�3F�u�w��� �%�O�� ����d�$�R�=u SN��q� �4��&���`�F�� \��M�zvT����(���	%Ѣ�|����R �=�_�9�] jl�㿓�4!��%\�p��`z�}W px۪E
3�xQ逝	�N�2 �F�Xڑ>� �h$�0������O���� )�%0~�!s�J`�g!cP���C�w K�&�:(��	�m^� �fy�S! �#cg�ܰ6q��\w� 
e���Q�@�a;�x &~.�k"P`� �>#�.q�*� U��R �a��@�O��F�4Y�� {�a6ml�t�C7����@���t�p�� )�K���QT�����L	@z����`@��O�wj����
��ڲ#+��;����.<Ϡ ���y|+8g��-��]}P�`i O��^eUh�N� �8��F
D�gdE��0��� �[���ch� �k, ��p�
��� �A�7� ��T`q� ��Z*� '�:2�rϊ����U��8�<>������$|��\Y�0�дw��P*��I	 m��F��M�� �"�n!��?�0���7{ �0�~���4��O�J�H�dd��A�?������q��@���\�j*U��b��R�0���{�
��h�9�!��I��h�=� �03gV�cy��д�-� m��<�G���l=K������W� 5�/��~e _0i�ۺ�A6���o����t�w��� ��̅�p�b 3�"���j��{ Uv�ew�Ջ�9��O�sn ж�]hG`�p�� N�sI�����f�����-�s*^ ׹�Y�U�� ���,2�<G�1b#��� �q��� ���Д�}>�@��tLJ�H(��`�x �R�TɁ��*W��D�:�$8�P��s `I�jղ� ��틓B0� ?J�l��G� 'yX�&����<��s��c� �_)ir��1�;�`\�0� �P��[�(����0�$��l��yv�fN�r=��0����> +f�6�i���pFB�V�> ���"u�N�|gl�q	�@�%��!w2ې� �eݼ�<Trf�O�^� l٣ [=}�b��=/f��DiF��S'W%I�@�!��
,��0 կǉ� +�u)<��Z �H*���[� �5����L����j�`u~ ]�f����� T��E�R�!0Q�Kk^ �tg��H� R;�}$~Sp��� _Y��ϗX��]���˺�� a�$b讃�"-�޶Q��mݴ �]�|x��th�& x�$���\Mh	��� ��B�R����֤f�x ^vb:����8 ��s�(/
� }��z��E��j�G�	є`9�Y/�0#�k �W�&� � -pXP�J1r���=	������F�RP,�ڟGx3r��27� �l<����L׾IP�X��F��e�"� �x�*<
d'����� �U7����,� q��=v��L;a�q[ ��SζЁ������z[tD��=F��6�����^� hI����}{&(<���F��?���y#�#4"�]� U.*�`]@Jp	o��n`t[�V�ȍC���ֺ�MZj��pxd�� �����z�=�z�����h( TK�@	3�y|����p���� �d��|ۯ �)xH��F���[���tHbZ�Ֆ�t i	��:�+, �ނ����� ��T��� O���cG�����(H� L��U큛��`2T@� ���n�����P؉�V�E cb���$��� "��]�{P nX��(� ��6i��I n�[���@����2K�.� �,;�v�]X�E����p4 �F��"~p# =eJ��7� �6f�����9�KVnL [y�Ǣ1�h̎�@"�>~	��t�@�j�nH@�Q�0�����;�@�rB��K؆� ��`�8_�� �@�g�q
 ����ޜ|�`}��t �,E(>�P��s���]�Q+ ��
ЦZ/�B����]0�_0w��ru	FÈ� �ϋ#�\�	}�:�X�M��(!�0��[ �L{�'⵸��T����[ �X]�G�Z=�	�_��W� \T��I�y�,�����힡�̍� ��(ú�p� ��*�Mz�_ ��K���( �@�N��Á �\;������ER��k �GjBғ�E >�Ɗ*�YAk�+ S�LH��; $'�l� ��W ޻F\�Ru��|�1��;�Z���_G ��nF���:o .�V�4�L� z��
���L5��"s�q��g�`B� }@�W
�� �iV��:���A尨P4�� �y�	� ��"Z2��E �6�V���K�
����v����ϴwU� ��^kN4�">� i�%0�F� ��GB2�� ;W�f!�|#�	�� �`V �@��HO������E�xr���d���&�| b�V���_�pW<�,�I MLw� t�c#U�p8�&���v.~9JrL� ���O7 A�*�D��㢍�'�a[��,J��Y��C��kĄ��������) ��p啕��m�밓"�4� =��1]�q��? �ƨ��8�{��h��I���A�M�Hƺ5 l'�m�W�� *��(�����f6�P �D�U����cB�? �1��P8�� ���i�K �+�W 0��^Ur .��lC��$�� ��/
��ٌ �_�� }���� ز{��?f '�JSbE�n" ��PT��*&@��$ x(y�7��l���5���t �A9ڤ�� g�.�X��`�4 ��D���l@`b ��P���Q B�o�c�] 䡬�C��2&/���"� �P �T�AQ�% �υ��+�&��)�_r�hsq�"� X=΀#����҈(��L1��8@�oc��&,:� ��lh� P`"&WM��?�8����4� �!��:d�7x�8x�1@�f�i�����
�$�Ť)Í�����TBt�`Հ)-���(� ���Ѣw+ ��u����1�=� Жh��, �R�ѻ�z� ��j	�	C��X x%9�� e.��| �3��M�9� Ѽ��rƚ� ⧱�p����(� �����L��0� ��@m(�2��J��H��<�}uP���u��teX��L�x��&�t�6.u�t �0-���|� [L��M ���VqE� ms��*~�:��u���p�nz�/���y8�|�~@`�vH qwB�ƥr2
���P���8����=4>[�Q�	n�p��ԔK�t2 ��Wq��J�=��V��ؗ|R57f��R�P]�֔M�3�ԯ���*{ ���p/ryx�wM)��� (gK�-���e�7:8�z�������ᤀ��� ��.?3��'������d��>� ��6����J <)�v��*r�P(\1$�(�Dw.P�B@�s��`��=Ȩs��vY�}�")�sa,��2!�A,�H|3T.~�<�!ceXu��:�	��R!s���$(�HT��IK��I��3�w�.�$��ay���(���� 0������
�$Y��`x9m[5
���@&�!��wV)�s�
|�>7�#ۯ�����\�n�B#'��+x�d��̗74��iܝ����D��%��x	i&�;  �Qّc��1 �he�a����}��? �г7 ��~�h&	[F�k@�4nh2@| ��@XxF5��H�O�h�uGT���?�t>`���H
HL�1#o�����������D��"�0&gN(�=qH�� �4ӯn�w�G����J�)���,�C4�g8��B���W0d8 ���F�Ek &��uv�T�&>�Ѐ6E.��: ��1�kd �SY(�wh� |�j��-n�5Q'@����} 6��ߵ����%�|��3���袳	�w^4|�@7h�v� �0�a߲By $��n�2`��@?<ۦT3� qU)Z�	bRz�N �*������9L�Z�2�� � ��1��m� �K�e��cU6�Y�`���nP� ���($�n��H��|x@0tc��ޑ`|��!	v �Z�"=h#��!����ށ1 a��@?���|bߝ{�]O��O�\:;��P�� ���PT���@M�����S� ��B �] ��M�-��' �`!~w?v�	sY����M�z�m��`�|�d ���_�n!oK�a�U; k5t��n�t1 ��m�u�I�J�� t��(]� d*m1"ǔ�H���G&��h��'����#5� dY������
��}v]������c�����I��"u���CH��Ӡ��� ޥ��Z��[�Ovn����m��PS �}�V�N 8�oXa���KuL��k�y@w����I�hޮ`�7 "�����O`� ��d���u�U�[ ����1#k,�F�e�݃���2�8�I\CQ� ��,`����uC j�o����z�-@���� F��ȇ�� �r�}ie!tsD�C��S��>w �_~A�	��0=
hH}$e�_����f� ��1�d���!E U��`�&7q���;X���G
p�A9�q!�p�vL��D�G C�Y�����(j�"'����i�0j�ZL	 A|��=1�{��B`0��HN>�#�LrpO�x�d@�ޜ�L��H,�� A�{1 :�%'�K� �,��J���x��� �a�u����Kr���5�| �	�_΂(� wHA6bx�`Lc=k�NB$qD �H&�1��tixէr�T	�8s��P�M�^����@��i��*��7���6}���@x�������%W��t�P�t�1~ݨC)� z�UAk��κ#8�m�	P�CLTti�x*Z���7�PE4`����iT`N%�f��~Ɂh6L�8-T2�h��P���o2��4(P� ��E7^��9�p?���&T���{C!��{��a0�1 ��Y�<P&\AT�����{:"���̞J[�im� �=H'H�?w *B��J�8��<��ش�/�t�i�E-H��y�T��]9��2 *�
C�;���,���%��ֆXC$��"��HQ&�� |@��4�����Ϝ��3	��pǹM0��y�U�T\� ����y�rp��Ԩ���*4�f< �J(��3�(XE��E��%�?y���- ��GS�6���`
H>��H5�p�'�N< fl=�"b6!�?���bh�jX���	�! ����|�(]t�<A9�#�Hw��������?� H8��&�KO��>!Q�|���e8�!��B��4�o �X���p�y�2��S�ƈ�$`�Y�I�9�4*W�!0Т}Bqp2�i��d��P� M>�����B2�;��^��*��:��) ��>8�R���5~���:y��0	��O�0>�Y�,�x��GLf�!d�>q`�);n� �
��2%	��	w��?*ǂ�|Bc�H�I!(���4�y$0�
v�X��O=2��0C� B��u��@I5�9�N9�ko�@6z?$�� �'�
�x����E� ���xvS��"L ��4@\=
�9�zs�2�ւ�5��:}Be{>	E#�j�υ���2C��4cM�< �}H|Ϲ�#<�1�C���@���	����O5��$? Z��۬(��;P�j�����2�L��+`�;�h��)�ۇ���E��c��P��u���I�u� �1�⎻���:C�7�!p���e�+CT�Ъ����nL"t",���@�F�W~��|0!LA��bY<�I���^ ��r=��Z� ��vӫPI�
�Ss��@4A �+�p6�T��s���`����Xэ]Ԭ�s��(5`b����Kт��8�ot_ e?VO��r� Di@L��J�}�ͺ� P��h���Z*����� �ɳ���P� Uq�lh#7> C����` �"����� _�~o|�/� )����E� 坍S���>������G� �=/���;�~��"}��ƀ�+��N]g��� r�jY��) [09by�۾z��	r�J|�����p���;	^3�!��� �HX�E����yk�h!`�8#i=8�q�]d�@�����-g��A?,p��J\�b���x���e�δ� |o�@z�����C8}Vx��TRLP�)q�L� :��{.�h��H�X9J pϦ 6fێdH�� M#C��q�{ a3�R�"ٴ �Ӫ�w�A ڿK�M��f 5rR��[ �צFâ����d��`ې�� �*]� �?�!��3Q��P�T��x$�Sn� �a�*�C0�M�����0:���tu� �3�����h`�)�l�[�}m��.	O� 4�� ��Da�(� A/E��0HW �^.����� )]:�4v�$0\�EF� ��_m�ӽ=��%uTx�n �(Z��N�Xa O���>0� �T����N0�Xo�] �nK-"|mb6���1��@�=��`�xͲRِ� �韨m�0l�h�T� U�`I8B�uC �ML���Y)^l�������� 'W�*�� b�Iy�d���/�>0n��#�":� ��wtʑ+��'� �4]��18�x�� �i!�<S�����F)�(��ȀJ�Z<0� e�Ϛ��x~���C�ր`�%�k�# ��LT9�/�B����,{UD�܃0 �E:\�!�< ��'�hTJ���1d�,�%.��(֧����i$��'�_��:Ž0> �yIM,�� �d^Œ�3P ]p�.��F&L�� ԰N=�z ����1E�b������;�:���H%(@��?����	=����q5P���o1��|�> ZW�EL� ��5y���)���H��Uh}`ɐ�k;�>:^#��7���E�0 ���U��;h��� �݀� ��佬�, �P��a�z����9�1��E���a�ĀN���� X��|��w� +b��7h��|�}�1@�����0=Y�)mD\� _��Q���b )�è���R j�Ъ�Ջ| *w�>��b��~�`�� $�>�Հ"���ӡ��tR�@pn���EAվ햴ޅ�0���kG�I�#v����i��uL��ɥ������j��B@�#�Wi���AqN��8X/T��"��H�$~<Y����4�F�Y 9���O~� �v�nR�]�m�� �x��X�qvր��pb���`�t2G D�z��c�1�� ƞ�(9 ����*x	�hR��4��1N�iG�����4�� p�UiCXD ����߻c�r��R���J �j��o��� 3�6:�DS �˞�	;�[����7���&q|: �5"'u� �KM�w�� �f�t�Z����@P���e�8/��1#'Q�JMd�}����̎��;�� F���e� D�H�K.pt��h��Z����LV��]0�`b�?M�cK@�p� X�+���`��I�@�>� �N�h\S{�Mq�4y��w���v [�ˇ�2jT��H L>
&�rD� �m.(�cw�Iį�5½�2 �N���ӛ� [(W���<S1 �m�]:y��p`�
R\�O����e%�� ��I�$|��d�� 7R檖L;��z�)�Х�u�	 �ʐ}c��<�
���p�N�wGn ���M`�xe��~�O��0k�2�����QchD\�6eX5jI )ѽf ���*�C�Y �Bq�nG�� ����ꍞ ��t��sO�O�&`��Fio 쇗n������"Nr��#��9\�� ʪ��m��x�}: �|H���ϢSbh�eq<�� ��V������*��=$��s�
ဨ֌�� �v��U3w�P��� ��ڎ�LL�tx U�7��} �g@T3�� ��K�tq Q$�0M �J�E��|G &��6��,� .b��2da� �D���	x������ �A�T\��;�� ɼ�I�X���c๳СE}<s��PZ������ ���w8�� ,i�+v���Q ��'����0 s�j��9A� �Ŕ�J��&U2��R� {��q��4�:m�����x`%1�d]�H�a�#ýR����Z��')f ��+R�F�g� �,�!� �wՙ����v�u�; P���ތ�����XV�$�]�d��r�H'?� ��6���p;8+�P[5.�=(m�� 8�4�� z.CPN���lp�n@�)�4 ea۱Udu� }H*�1��-�L��d�:�ǁpqjk��Y�V���5RCK�U�:{�8|�}'�iu��Mc�v���Р،��-u�R_m`�%c돰@��/� �t�?���p �l��� Y�}�76� ��&�%�� .��}_�/��z��!*�^(���%T#�� ����' ��T>�����f�^�@#+��b�S�,��@��� ���F)$ \�#��rO�nP?��GĀ(�A��S���wZ� �TV$z7E���b�/f^�R�:=�� g�nV���+ urH3}� �*��;� �:�Bfì� Q%��v��^˰��������y� ҽ.<���>J����| &��,}7*R?~q�#�|�e��yz�Lb�3���(J0<� ����#e��(��� ��ڵ��g4 ��#�l�G�H2��X���@Ɛ� \�M/��4��@��U]� 0�	��� �i9)_�2
ӚЮ���:��딜���Gw�<U� ��K(� 7jaCY�8���v%����u ۵��τ޲ �³�	���ˋ���}#f[��-b �����4<+(�>$ r���� �N�=��~�W;'Y Ɂ`�y������K� Z`�<t�l��_S^��u0 ������~� l��>��P��]%E�?����1-[���8�� ��D���� Խ���jF'H���@w1A�|�����C ���6�x !�%I� DFA ���ݸ� ��X�|�9���ӵ`��B�E�����Ȟ�8 0����Uзb����+���^��:�#�����|�7�F<zMX4 �UJ>�}������ � �P��+S ��r��%��e@�{��P �}���\S� Z�	�s����� 
)�!(� ��T��@��H�� 3�h��HǙ�� 
�^8 W�q�(l˾��$�x
y'�-����sָ��V o>�6��B���a�0�M� �TJoI� |صXŜ� �
"��h, ��5�[�x Zq���ct��0�J�်!@��yt� x�:5��� ���z���� A,��9�.� ��y����)
~H���� ���_��p ��EH�� ���s��� F�-0�i �x����}@)�����`�, ��{��6(湜��$s��܃#��� �&U�h  I�S}�D �@��H��A%�&G���or����Вb� t"*�8��^�����Ľ=xX|�����Фd��C���l�� �jnXwg0��bo�ؠ0�p�q�P#��}�%� 2�x���6��9UW��~����� ��?' w�5.�!�s]N�R�g���p��;)��	��\�����h� 4�}[�Zy�P;r
�v�����T*
� �<lj5��| ��s�F�!HEQ���,��� �I���k�y �׋)�-� ���vU��щ?�C	�_@t�_�) ��~N�]4��50�n�'�7`p�9����E@�i�ɿڐ����p���,��̈́U �Q���G '�F�YX� A.t�(� ��V��W^�MGH ���.�q�{� Ʈ�~�����mh�<p }��ǃ��@�?� �ʱ�[U� �5�T��Qf��m�����)�o=X����]e�Bi �A���g7JY�[�0��@�3�S��RW8���߉��� ��a"� +1#jY�� �SV��?A.�~� �F�b+��� �8�rc���w dI�S�\T��U��M�9 #�	6��;����!}�4E��ߐb��Lu� r�,��(F ���a��q`3p���	#��F�!�*��Є�����wg�Y	N���U�[�)F��yP<�� qzc�N �d���t �b�y>?�C8�����B�vD��9,�}��=�ـ�鞣JtW�o��O�)�L "��/��>�.�h��WƠ �~�f�#pU���eyg�] b���(J� H�:ݏW��~d�� �
%�B^ {�T�c��� ]�A�� �h56@�`�`����s�D���sB�M�b������ A��k]�ؖC����I���f	zP�e��ĳ
��x�8~�`N� ���X�o� Kƀ\��]�C�߇`�Da�ѩ!R �d�'R8�b#��A�V����G ��ą�X^��_�A� ͬ$r��k�  �ĵ��� xe2��|* vѨ3V:/;X����@���Y �^
�S��!�@$�W�s} �y.�Bn�D ��x<��0 7ȩ�N];?\��Dl�k��������_�C�0&O(��y �ǎ��'+� �T;������
��O�+e8�P-0|<��0�X�,q1 +���%�6 0�ә7�w9��aN ��`f��<z2 ՠ�!_Cr������"i̶�7aJ:02e=� �'�p� �I�"�E�l-R�g7��7b�`����mH��{ah�4�b��ҩ����6��
������BZ~�:˩DԾ� C�m��7� �����H ]����#� �$�8
�;n�@�[핢u!R���q_1� s��� �gF�Q���
q��P����Bs01r�����2��4vЇ�M� ����lF� g�}q�?% �'�~�
�. ts��oC �3�/!�~<�J��Vg���C^f������
��	Ê�)5�b�����J�ÞG�QLD�A2��(r!,@g0D��0�x����b�c �k�x�1��)ڛ�w�y�j)D�.ncy�v)܆ �1B�QK����D)Jv��t��B	�*� ���h�0�_���K廀�Ӱe6C	����R` n�ۅ�7�Y`G<)c�F
l]�p� �;���+K6����� ������Ut�㡛��L ��К��� <�Q��E�r b/20H#'� �WA��|��!� ���9$l���� %b��7 �&���m ��E$Ҹ�9+� �- ^��p�(M5�����q ����v)�{	 9ɹ]��� ����c����qu��a��� mC
���	&��*�?V�� Df�e���;h�
��|!�� >�=+��G ~[Ү���� �h������ ?�`T�� 8��0Q?ݥ �.:����9�ր�R�F5� '����-3�I �
u���1 ˱m�c�D ���
8NB 9`z�}?;��L],�l	 r{�<��z6 +Fߐ�飥 �����y��0@A�� �SU�kN�y
�O ��s�G{�<��)�] �� d��W�����S�����?�� ���L�8��wg #����/� bX���W@�8j��F���`:�Y�J���I� 3�b��>�. �?�{�RJ ebg�p�� �����R� ���b������1
S)~%9�# gh��K���QMR�q� 
F5c8p* ͐��ϯ�p� .܂�� [՝���P��@�:
�i�h�3��� m]>��Iw�g<0Ċ�X��p�"�Dˏ ahk?���  �UK�g �Cd�W�~ ��%ܥ	]�-��@D �� ��7Zj�� U���Q��, �Ic�%H A2�d�v� 9Žiu|�"kO�^+W@�=���&D�A@;���@�N�<U]�S���-[6 ��YC�N��x���� �)�,}�Bu� ����H �6
��� e$��-N4ؿ��а��� U��uv-�~��@|��(r�y8 qAl�ϔ� ԟh�(_	P��3���R���`x� �u���9�� 0p	ƀ�1 ���a�L�{� ���\��v�y� -j��r�ƒ��^X��Z=� Źv� ��yI`:�J_%A�� d� ��["��� ����C`���������4.�&v�H"������ � g$�,�����\{� ������BP� �X���j��J׏�����te �a|�>{P �)(� "�_����Y �b��l +�A6ˁ�z����&@�"7ne�F�.GJ�@R6�\&� ^��� Ϋm"#ϖ��� i0V�k� -a�P��c����s��g p� X�{F^�( p�s�'� q09�a�^ (c�rn �וHv�\�˳����n	\� �s�(Pe�S	h�� 0�W� ��(�M�
> �8���{:1�����pW�ȸ�Pbvbs� M� ��x�������sTyq�jX�@�P% ��<�on$� v�8_�p� /b�Hw� U�:S|��� �i���EBLF@;8�q��_��/)`"�i9 '���f��PM�ǵ 3q��[8� ����������I��)ڍ� �o.�Xҗ� �}\���I �!hU���q��� c�l)��F��`Iz���&|�t K�1x� �L��҂mB <���c�xQ�I����ױ>,����L����<�%L� ��g��$F��x 6�v��&���@A�{e!*u��M���b �a����kD���ipAC<@+����{�w,@������&xG#
�`��t�:�9�i͎�88�� �����*�x �w_ׇG�}7��9Z D=�6�1PE������Q���I���ݦ��d ��k��s�	p�nߎ��a�p)��#�%��Ҍߦ���] �r��ʾy �h2L�w�:�� i��+z�-g�a���\%��Z�iWP��� ���o�</wݶ�'r���2`$]+��g�������	�d�� Z7��g�& _z��i�� u ���a� \��,� �mtT�Y�z ��q��Lw ��	�a�1e.ǥj{��<�� ^�9s�ģ�u"�� jb�g1X;>o� yAt�T~XP Ħ3(� !��ݖc� ˥��o|�`<æQ�MkL� 4�����O7 Jq��]tX�� l�o�*Z���@v7 �W�?rm0� (��w�8��� m��2I �&����q� �ia"�2�B�}� EeR�-�7t����W����1p�V���I+�����- |U����}�i�� J���`g<�tGH$�9���q�A`_W28� �TV"�=�H�`Ol���1 P��8y6�{L!$��~-@�ji %��l�, J�� ��0�ܮ�O�����]� ���%`�Ld` �;A0f 37M�o��4��l,����r��=j�\�*�>�dE�(J�N��S�D�� n���L������0$?���N&H���} ө���y0�EPP���s�Z'����c�W[�y2���\j/��� �.�n��d3�`�[�z� ��0��G̪#��s�4� �U����S` �	�+:�V K����j [��;�6���E�����	��� 	�x g2����� �;m1��-9րE��P�����@%e`��=�= �D��X^C *h�잕{fybcMĀJQ��� R��UT�2�ݎ�W\B) ���iD�9�Ͽl �?�պ��o��,���)�|� R�bCD�{$ >	BG��u�*�!��6 c���m���]��@��`d�"� sZ�|�Ϣ�0�=��P��� �"u�qH��#d]��Iv�HX� � 4�������^�w7�` ����3 d�C� 	�V L_,��*�xo ���ԇ�G��EVI/���Sx�� 0%�Zd�y� ��H�f9� &a<}5��7 �1p���l[�~z@
Z�6̽F��� 2�$�q�V �N�p�k ��;���:� �٭���S*.q���R  l�y�$#��������w�Y���cb��k� �@�������R8eЧ�yn��B`�[�P� ��G=,�� ���"��� �MӡPZ\1;苀JΤ��/	"��	SR��@�9Z3U��8S�V��wv ���17� o[��f��>�&��pmQ�`j����} ?W���p ����Q-��b;V̂�Uj��@�.�`y��J�{U���bf�p`�!E��3l@�-�똈{���'p�`��\��ǋWsI��h� �eї�"���8,���� �&�>Ӟ�  'Ik��Ƨ8iK襲T ���Ѹ� E�9-&	���y�P�!�� ���T�(9 ��/b�� Oqi��T �Ύ/x  �p}̝�D�2��g? �F�帢a��U�p�tM �E�r��� �H�S\�N&C��������n?,��0c�F s��woq<�6 @�IʉJ�X!pF�{�� ��%aCw� M�H�`�[ O����>c� %��K�=�*1� �?9�NvG;K� �c�-* a)vI��� � >"ύ�� #ց噄H �0�pu/+&&��  �f�8J~&0o %�"A1HwF r���� �X����x���G�wFh��J�Lkc��'xF�dc���ĝ0s����L»`%�(����P0�f� S�O=C՝ ���ܳ� Q׀�z���p�Rij�I@�Sy' �[�~OV��Х�}����6p]`�� �PU�y Ӫ�2?msI��ڀ_�r�ţ����R��L�z�
[��t� �싼��\���k�>��3�+0�#���: ��*F8s�� %�1I`
� Z]�HW	��5�@�� ೈ[�]��� �7(ڸ�>�ǔÐ'w<'O��r���	�f�'��]���0� �𡺶�3� �m��N�� L�~� _�;�y1�b ��Z5� �j7�D=B� �G����D�,�0�m ܘ@X�i (J�T������<R �֥� �AJ���t��)�J�G���0��*�>�!�a@&�U��ES ����" q J_�������Gj1��vJ�`H� P%u��[� Ұm��2$s�0�ꠐ�Vߺ#wu�x �mB�]�.�Ï6Oy��q ���4�br ځIgT�0x~	�&Ӯ����P?�a �ˣ��L C����� ����fN [�'yL�{$ +���g�� ��h�� ��T�O�� ,�t��E  ���6!� d�����]. ��2��{�*���$���p|R��<�1���}����������Ͽh�ة3�ףB ���%85D���	�� 
�����'�����jm� k�V�	Xy� |+.�@F�u�Py; cH_�G� �(����?Р��� ����Mc� >��\��]�2`r��� +��ŋWs� �a�� �$��M
 1�8喧��R���@��wڞ�_��8 ��3�:� J����� �M��I3 Oo��Q`;�� ��� q�$��
	X�q	��πp��� �AO+��M�N8^� `$��\��� �'�aɰ( �攵�;�U�-P2�� ^5��Y���X���s�. �oߎ�в� $4�b�{� �
���� 2BrF���������_h@ ��&�*� ����5�A��h�(,y�����p�QJ�׀s�\Č:�[�(��l� ������N��{�< T����l���9.%�Q�H
 Z�}�cp�=�(�$��&�F$@-�թ:�,������h
 ��vk?x� �;X�,��]Q�̐�9R� �I����[f�i�nE� ��X�	�XM�D��Uc?d�
��~�� �ˀ=�!_=� �(0�L <�k��
 ��8r2c.�$m �Ԑ� 	��/ ��?� ��hșkV�N|�����`�(�xX �e��O� �n��l#uD������`� R-���ې�wJ	���DHx PCF%�<�]�5�A}�����)��#N�� fͥ9x\J�@A�U� �ǁO�&3� ���f�bT��,�@���W����c�zlm��^ [�{J�|W �˝��8�=`4]6���E8�)u ���(o 
f����|� |��ag<�� !F��9��B*r; r��:�/ ��8#A}� �X�d��� �SB��px; �N�R�=X 3* ��`��@�ے(M �=e�����)��3�lԀ�ZF�� ���UB� !,��#^�X�s���}�e�����d�cհu&� $��y:�tR Ow� �-�~8E��$���?؊*@��Q# �'"t.?�sz� }�x~q�j,�[ g���J��y���vP�4p��V�_-�M��
x �~rd�cs #��+q�� �F���w� #�שZ ��.y'���t�!f��o�r �k�L��} ؉��,�՛"&�v��ܟu�U^_�p`(6-�7�'��o���w|�	�v� ��	u �M�W�S� $�pV�bKk N�F� Ct�x�蘨���;�bD E����<�z�L��g����̤F $ ���4�{��pc�=�- ����j��r� w�Q�.U Ng�=�^�{���s�,a �9���A�����X:�d�-�ܥp���t�"�(S;�� y��7+��XǕ �*ҡ��� ��a�>� �t���8�� �#Ybn/M;�8�B�@�2�+rAC��/�?o� �WY�RO���� �	<�1Y�\��e,"(`�"�� �p�X}��yŮ�E���5 j8�)��:�Q�(fT��u��3@��Y��	�&� L��U��u� Z���el�� sP{^���C+��b�r@ $���y �;]%v�0 䫈O� m����M&���w�V��DG:��u��= ��/$�� �pc�o�(���V��hT�� ���#��� �Z�A�L���Q&����'C���L�P$fV�Y;Ѕ�� �IRPϕ 9q4���(L�� �R��}��� ��̪e1~ ���ٖZ ݨ �zR px����� ����1��bL/��$�8�q@�tT� ��6.P���z/�L'���� d:
\띀I`#O N���.� �Y��>���0v�by� ���T��=��!S� �aK�m{
�� ��}V��9 ��y��~����AB��\� ��ʘI;�� Ɉ���
T� ���3�q ��:�0�� 2j�/��\\*Zy ��4u� �P�tgֳ�T l�����b #$�=��\�MO��.$��Ȁ-RmT/ �x��;\�*	�B,| �^�Rc�!����H)���dY� J��G5u�ÖV�8 ���=���8��U������ c�!���^� l�5�xz ����{� �'-��)�<8���bG��f�6�r�0@�]�����=�����q[ ��#c�
�,��� Y���� 6���A\ ٥1���� �0�@Cd�W�� o!��� ,E=O0Z^% ��X�ia� �H����+� ��«�$Z�> ��ː�F��<1���� 4������ +;���?0vKD�A QJ����Iq5 ,y�$�; �l짔�� ja�<C�� .���9Y~y�ܨ�@][�+�����)��m"׌�+ �'��	 �#��4�9J �E��S��p͜}�Ѫ�Ƚ2���QE��pW/Ѳ7�I�'{t����� �w��� ��Ik�SP~ ��j��˓�� Yy�(�Kd2O��h�٫N��V Iz�H�v� x���!�� �D�sT��� ���h�@� ׹E�� _���u�DH��zN�� (P�:��" u���~�B ;췪�U�
 jL�tg�=�t���k� ����;���8� {At��̀��RV ��$;���� �O���^<�� d�t���o�r�� C�0�Y��Uz �'h�9~-G����L�� ��0:d�	��k�Ш �2q�X+rvoLw���WH�s�q���
�� ��R%�隀GY��]� �*����Eq�f�9kܷN,*xT���� ��Hu]�>�9��>�a�|�2���b���:�[a�	�rx� ��^ig��� o��$�� �\� H���<��?�f=m�	���� \L�;����ꈰ̅z��M�5����F�DWr�i��h U��G:�I ����k�� ?T'u����\��%�`��b����G�+^P|v� "�e��D= ��>?_�s8	�T� �U�4 ��DA	%� 
�]`M�J�	KE�8�7 ��cJLsH�p ܷ�{�8�ۀU�#�?�M��/A�
Ш��� +b@� _ ,$Y�����CV��� � �KP��EFb ѕ~q��Q �<����O%5��vZ��2O��l�r t�c�=JqA�� 㨎�v� eګ`����HGa �{��� ��<���� ��E�0���G.�(� ��񢪼�# ��V��iYyR	.��ؘ 0���䍛� �~,�<��8���C�`�'�32��[� �u|� /mM	l�
�n� %*oz� �b�ӹ�����g�>}���}�2^���O�ę����M�#G{3��q�����]�'P%<W����9 4:;1 {Z����G��fyF k��̾�� �+�LO YVF��M^� &���	L�A�3�p �����!�\_�r�^����wK�(�;�R�r�����wB�f`L�$�:��b���*�׃���二�����מգ���}>����YZ��hTE�N; ���N���b�aI�vjb}�g�H��!L߅ ���:#�I�C��~ 溝���w����� �l3�ۅ� S85+Tb���1o�t�J	̜��TXV�� #H�'��C�0�"J;
c6޿���& ݝ"�D��°�
}�%p��8�����Vx;���R� �� ��?�(��>	X`�U����J+	ΙE=���b��o��_�� >����7� %��:��+X h$�x4� �_J.9wc ��gۘ� 0$�8�q -�W?#���a @�GΡ\
� v3R�C��g�	 ��Ə�Bqdķ� ���ŝ�;\�� ʉ��#�"��w��c�z�١�����ܛ ����K�� �(U|ֻ�	8o� ��B~i ��VO3x*� �#��H�;�dW�A��> �7�[8���X��J�D�ZXo��[@�n^� ��!�/C, @j��A{+	�6 ���x�V� k K������J �����v� �_'��%V r�j��9Ju�>�R���B�M��@�1��gt ެ%j��] CD��&��\F� �yt�T��4؎(1���QW�h �g����)czF�_���K~|��%��V��?� Tf!��vb� �<?=Y��� ���: نfˉ2���� �aݸ�C Ml�F��+A$&�ft�Ƈ� 7�jl�� �=�;m{�s ��t���_n�~�� CoN�DE� ��B���J���P$ا ��"�In �/���o��>�8 ġ�d��.�(�'��	F�LV��@�3� ������1	n�o��@x�~�D�)S ��<dٿ: u�۩ژYp����Q���~ Pu�co��"mJ{��^�O� ��`��,��@�.� شZy`C�� �W6v=��� n�,�.BM\���� ���@�� � �'C�_�.����vi���� M6w8ة�P�,;V�Sc� /<�Tô� Hq?N�*P��` r�s��h�,�FbcY*��Ѝ� [�ІpU�3mP�.�֬��BZq]��o�L���)��� ^��{�Ħ� 9����k�b L�����_ �1,��eG�+(2༤��� �'���8T�|\V�"X� y S%���cӁ�-2����)� ��h�D� �u����a~y+��@�ȕ���� �4�R�r�$'�iuLj��z �l��v 7��m>Nu��a����,2�\ ־�
�ƩO ��j>�d�� D���$��H�9��� �<����% �.�3O"� Fqϰ�?`��� �T"��vX8���� �G� b�|�7�) ז�X�`(����L~<�p	P!z c��O0���YR^�Ǎ�k~��y�+B���آT���4 V���l�m_�
@`8��pC�} �|�h��*$r>��5g Թ��6�9�(���-�!�� �����NrS�ʛ� �����	��0�Q �-J���8�Ԃם6���.��A� �]b�9=�� G6�.KS� ���)��uo ��m�� \��Nln$	�� �P鴚{� �\s>,߈� ���c��e;尀&2��^�|��EĠ����� ����\�	���� p���#	�I- ���� ����8	� ��
j\���5 xB����SQrkFD�� !G�.����Q�; =�d��� I�m��t$�kY]�poU�*�� hx/K��| �ϵ�#ܑ� ߁Ιۈ�q �Y_�Dz����ᐯ���̤����Ƀ�@�_�@uL�k b����h�~� �}�O�d� �F�C&����9��E�U� �O;1'h�-N���qZx���V1�+�]�09-5��^��� 6���qW:*C���T$�=}�_��J0�^4��b
+�� U'�T3��j4]���K� u�GJ���; ���,�%�4�_�u���jH�� �&c�[�":�j`�§ Cȿ�m��F�?���H��� ��K_l�0�Mk�D苒� ��T�y�	�O�� ����/ v&�^Q��`�A ��+[}�Jr�Q	�4 <�n|zր ��ͅ5H $��lF� <\�����L�~ #�!�%}v�������I�@� ��D:7�(��;T�M��=% *��i_ː�~m4�p�&q�Q ���%�-�e�c '����ly�h�1�%Į�8��L��!Q���g�vI�]K� }����fL ~VQ�k&	(�D(x�8�@������q �E��XhGS:�]��^�1���Y� sm�$��Ix4up��~n�=���Zأ�� �,E2��$ 縖J��DvV�u�Z�� �	WnL� ӦRx�т��A����n@Rsܬ� ��g�� y*�ѥ�"N=瀯��f�D��v
� �T���&��/� ��'��� -	�0,�� S���#Qݹ��p���V �$THi��	R��� �ܘ#� N�
�no`�_>yp&s� �M&�4� �ѣ���� ������ >���4���0�5A�mr|��. ��ό0� ]������=u��5`堌�cMP�|�NxaWv����.���wS p�|�׍֐��3��(]�ha у��[X+ lxKG�Q�� ����Z� �`"8y�� �	j�4Dn&��l�G��� �W�A�&zm���R, w�M2�� m(��Π���/Ӫ#��8; ����9��e��'�z�r�6������
��� �2�	� 9�ņB+���zp��W*��YK�HN��x<�>�����(ER[A ��s���`� 5iB��) >S�@$� va��C	 ���l��0A �v��?+� O^*9�3���l�S `�-,����Sqˠm�tG?��,�y��qg� >�w4�`�? �F��r��� ������� �i�k�Mb@;՟��{�E����;\��"Q�7	0�� �w� �\�_9� L7����gtm�h�Xi���$����4ܖ '���R` ��fd����5 �՜�L�4�Y��Fʩ�^�M�&lg! �����,@dа�W h����~ �D��@Υ��9%p��0�� f��W�>S���6�u���1]-�	��c o'H�;~�n2{���wV �I<� S^�C딀f�qM�t� �Ya�·�$�ɞC�_�e ���#Xg)1��Ӡ� ����	�d6�{��}��>��: �d��C��$�6� L}��.�[򀾃v�;od������Ѱ�׎��X�F8e�0�H �vcTĮR	 �59x��pYy�^PR؂� gdC���� �[��W��L�3��	z��:- �t��[mJ��>jW>�<b�E�g�LcY ǲ<,M. �`%l���)�9��ꁞ\:o���pg�UB���X�?��`�jt�S�d�� �}����r������`�N)o�����Y*�@���rbĄ� �U��d��� y@�ZB�� �CKp���i ]�%yR �l��W�I$ ��=;ɁN�y à��E� '2�!���t?����Mhu�*��	���|�\� ������!p]����F��E*���8��8Y������W$ ��~��=g>-} ��'�!n;�qZk�`�۠�ً8O,�� �9��� ]� k�K^<���Q���+� �O�®�^ ksh�=1�y� �)�CƘO }����-�mQ��d���d�v�_a��@-0 �,6R�\�o�}�� ,����Ҳ�`���XE��䀍�$�`?9� ��S6����H�aP˭�Q F�޴BC&fi�� 4b�Q� 	Α��9�ԋ�;���k��=�ȑ�{�<�!��x�̣����f�M��hB$��@A5ۑ�[ ��	����D" �yɄ�} u�VUL�I�~x ���_\��^nԤ'7#��&�0�,ja z~��Sv5 �jb ��ͷ�8�� �X�r�H>�t��Ka����([T�@�`�������/גb��a\��� $� ��qi�x�Zt�}=E �*�> ñ�W�m�	�o�D�Y�0�؈���0���|H v���G�3$�io �^�U�7tf �x0�n� ��V������H��@$�� $��I�N K�#9é�� �+�Y]����5@Fo�D�±����M�W�2�[R�"6Cj��fI`�*x� BO��X!�q �M2�A� fT�[b��|��rFuo�֪ ;=�m��� M7�����i⠼�+�:(�)��?�G�<��8�3�p� ����H��������H` �<�4RX�l(�����n{� TXOC�J=,� ��9*��~ �o=myH� ),�^f�{�? ��/|Yw� C�(�h�H� I]Ö���� �G%�0W�C�g� M���9��r�!K\O �3^Tw7� b2���`$ �Luo�@ ���I� �k#]V*����@����yi =�ܵ��� �J~,M|U y�^��P�	��� �螦 l-�6h�:ܫO�a��n����#u] sS�1B!�xT9��D7�{���>� ġ�� ��B2��L�� �h�]��� �D�k��>� ��W�9 ���nN%j ����� 7R��̽i� ^��kt�, �:�P������bW�;:j�>����0���]��ơ��0���� ���4C^�g`� 5ݍ_0��
 �(���}^xO���>�Ф�I�;�� D^�?����Xǐ��-� �CQ ;! ?ZA���$}`q@D��һ R5�hs�\��_v1��}�I �&�Z�� ���;��jD%���G@t� )���J� �E�6��A
��Fcȇ?@ |�V�s�� ��kA�� qFN@58H_L�
���8���o���I�	� ��86 @�o�s�WHi� ��v��P �p@(�0�� �r#�b�� �u���(�z=�1�'� :H0��s��>�W4�8؁M �?�ҝ��*�� �4�� ��	�X����y�Ma��@��(c P`W6�),��� ���o%��V� f���?���簈L�Xc� ēTd J�䍒@1�� ?�[ڗ��� 0G�9+=�����p����5��_Z ��=�i�ux�;9�ãÅ���`@�Pg( d�=WǇ9#n��-K����&�x�x�s�cθ߬�ـy`K^ ��\�L�%�A�l]� �$B������^!�Ydi�g�L� Ĵ���t�[ q��a��) ����C��O`RY�%�y �rk��� vB)�(_ ڥ��r��q p����.� �Y�5�Q�q�O|��P�0�`�A�x�5���eH��QI� �\�;n��XR���H�Q�ې@��0&�Ș:Ж��� ��H��ԓz� G-�Q>�]����U �8���n��aq�O<_���� 9�^��hG�'���� ��$�晈<k�Zqa�� $��-��b� ��$V� hN�U��C q8b���=?Ä�E����Z����P� .T�3�)$�TY�+� �����.L d�"&zl_u ө�SNY@ >����? �|GUT���=#���z!Ds��̏�r3��͢ ��8�Y����$׹�OAC"V�r�Bb9nT#��*K �}N0�u�c��D� �F�d�5H`
���8�jK2x �.�lKF��H p�k��\�1 H��B� ��T:$��-�.yӟ�����s �,X��S�T�) 3�����gl$�9J=��e�mQ�|�A� 4��p��� �T�1��`$"� �J�k�h �����?a��S���J`�񠻃%�� ��Y�n
��o{D�P��t^	M?V� ?'�� bX�9�vZm �;ҖH�h �ღ�o� �1����}G�ݠ%�\�� �徛�4a<�m�6��Ň�%�� j��.V�?�v�D�� �U#�L ����t���� �O��7�[1�0��1��!��?��o l}��t �hC��w ��I�	�:Y��É�d0ZHXNu�o��2� ؉�� ��3m~�>xe�Q����P�ճ�� � �(�Li��=ş���� �\��� F�+ozd�e��b@�<�(��� ����'��j �R��U�i�\P� o	�}폂 �xT�!�~d;��Ii�8����V��K�Nuw a�	7
yb fW�4��]u H�v�ӤQe �AD�Ԧ���\�]w�Μ~�(��^�z��a��Vو\����)�Y�b ��~�U� Skg��� 1u��m ~rډe7��[ �9]:� pƧ@�t� 3u�J��y� �qⱂ�i\^U�b	-}���#} 3�4܏�~� |�ۑ��W�(�ED<�HxAO��N�(���t���[� -�+Y��)e<�b�
���m/��\��,�� ��ci�Ƌ�������&'y� >	
��Qra ��E8;d�  ���p��� ��O3� �����9y� XeT8�g�^q�$]�� (��� �h���IQ y��M�����р��KO^ ȷH�&�� b��:���
 ���P�y=��.I�j� aC,^g	}'�hM���訕	�|���C��g�-z~�!��+x�հ��@�e �����&<Lp�K���4R ��'-~L�K@�l��� N6�O�o� ��fu��� VCt��y&,OW ��G�~Bg��܀����) ��T�� ��<���^ �7:�k~C��,��� ����� rQt��(� �2��vs��@�RҀ�E'�� �����]D	���}
���� |���#��	�
�� ���A��j3ϐuY	� ��T�Z�S� �����I b�M+|�u��xGQ��8v�{c^��\�b�����UK`݌�� y#礎�!�_f�B�$���9����/���M)vQ�$g�:��H� j���"�� �`�ϙ�U�� ����=?Ẁ��#5��] T� È��� iE*��[� uqׁ��y�4��& I�F�.v�O �n�$}4 ��#���� ����PkEb}@+sT�%�[�����mf� �~�I��UV,]�� r�"! ����j# �? k�a�q ɻ��0���$p�6T�uoj�( &��?�Xx�؈�^ �HC�P�����#���O@ ���݊��F�me`�"PT� �u�6��0�Ĳ"X�����H�� <�����z��x�0�W� ���Y� C��;X�� B>�z)� E6�����rI�6f=Q�_1�~�W� �8���$d� �(q
�LA���,�6ף��g ��;��"�~�	i���+� � g���2� GsFV�� jM�K���� 럡��f( �VE��9�=^~T:u�`ٍ���Àh_"���J�I��0�
�T O\�5W� ��i�D��$�l� 
7����	h�� +��٫�A5yj���� ^�+u_�<;a�U:����s$������51��Ӏ
�� !x��b���F�	@C#�IN�5۳��A؍?�G��i��t��|� ��[Ƈg��~}� Uaq7�)� �\��N� z�B6�j�� �K��w~� |\-�oH0Č���@��U ��T3
ﵔw� wz��'��% t�:�Ԟ���6u"��2{� ��R� c�S�ר	i	B��\�Y��ݴ E�0+{����I-�@�1�z� ��Y(�ؠ �dZ�!��� �s/�lX� ����Y m���c�� ��{��n�A(����=>�!X\���zBV��@�y �Й��Y ��d��7�(ۥG��C�u�0 �N���L�|nQ��Ȁ-��p1���,�� ag�eG�"~�%!MT�\�S ���@��H�-n�x 9��Ƒ ���tH���&�1#�� �}���m3A�o�����B{`��
%H��&���\s<5���3y�#C{ �hg����� X���qR0�p ݽI ��HtB� Ġ�E�n�/ M�
h��N)��������?�D�O<��l�=9�1M��e �q�"+.�� s���!/x�&��� H�uz��X�� 0��r���<���(z*�/9j� �+����a2��L��p� ���%\�& ݬ�?�Z������>����I�M 6Ր�貋<��Q����6�q x#oz�gw}  ������ W��{J��( ����hXv NY�+c�E ߬7��Z|����)G��� �@�&wƴF�b/��"΂DL>l��6�H���D�O�Q������������ R^៘��K ��5�H+w��|���?��~ �W����_,U�c;&�� ȕ�Ϸ� ^��$�)Z ��r	��Af?V[�X���7 �a�ޟн������ �Pm� n5��ෟ� N(���yT��p��z �u�,� ��C&Gj+�0���10K&m@ 2a�U�;���T}��l �����i~�� sfOޗ}�l~{M�;���� �e�� N�vѾ�g� |�
��K������/ܝ �SGz�v�L%��o�Cз�7�	W�dwx ��(j	[�0f\c�"N�Q|�I?ǲ9�p�k�� <��� _e���`� HU�r� �7��exL ۘ�$��n {��;�٬^7/��x�R`�y��8�W�� \/����n�1����H���.��-�T��@7���];v �q�Yo��� 9��P�� �t��(ә��z��V��t6�i�� ������{ ���P��ю�
e �4x�X�8�n$7t�u���Ls�eEY���\Z����� �߽=���� )<@�w� �1�	^3����V>͍�i5`���Ng���A��b�4Y �<�G$R] ����6��U<ܠ� k�4��̲� 죚n�۽*Q#��:��U�K ࣠@  ���k�hlL8�o��]t Z2�� �}Y�����
O �-��m ���s��� ��6l�p0D)��� s��>����� ��&
0� �'�;@ ��S���QP 5�qk�&�' u���O(W93� �<���	Xʗ����hx��gdW��lE m�+��M�o UH�[P>_i1�zw k�#��?�
���A9�z�n@���<�X=���A� �k?��.�� �T
��� $�����LXK<� l�\-i9b���)q����W�^�# ��0�s� 7f6�F���r� �ݹ�V��-6���^�頸�t�HϺ� TK�{ ��쁸�� w�h��U�H [ț	N��u|�)������1��UӜ ��R;-�� H��i���y?6�zTԀ�I�q�b)֮����G{?w-��a �@[���G��X�* ��T?iy���u�\�!�W$r�b�~J��q8���E4�m�
��tPc�k0~4������� �&���,e�` ���?t TB���A�J���`0� �H�'n������ �l�N���Ekĉ����Swq�T@��s�m �o�(F� ���|ę����ƃ���Vg )NnP�! ��/-��� ^�ړɡ#�;�_�M�.h� ��~H��%� m�.�,�� ��i��� �6��U�>ӻ�� �y ��Х ���r��� �@�ա�hp�����MƠD�� ��<(��� �'.��9}� �ЂTf<� Ϯ^I�$1c g����M�� BK����� D���t��Es��o�%|�  �̋�0Z� �+���y�>��ih �N	 �a�6�X���B�|��p�ݐ�� ��ɖ�Y �'WZ΃_i���� z����3 9��(>B�����26�eH���y���*9���W ����JU�� Y�H����ҭ��S��_q�[�Y@��k{)�~u��;�0# �3xwEn �ւ����m�OR��ӛ��r� ���!�"�, �9�)�� �|�n�m��y�G[bu�p	I�  }��7d��6 [Y��� ���R�Dz�p����F�}E�7e@$V"mr�a⥋�}y�9�jis������Vy� �>N�&&ԥ�ເ.(ژ�L�� @l�g��� �p���c0� ���ԅ�SF n�<X���W ���&q�� -�� ]�u� ��_`S{V0d�֞�b�Mj���� +Z�T��"��0��R ݡ3��� ��w�1L� lY��gH{'Aŀ�k�M3�� �<��Lշ&�:x��]�@� hN�sv֋ '*��D�R���
)E�L� ���z4w�C6`'�O��E���Wj���-l�`����A �1�t�v]�.� l���� �@#B�V	M�� �����,��t�E��D�<�W �x����<ὀ�y|�&�� �~��Q�� S�Z���(� >�z�EF%� ��逬�.wf�!�D���?~0 �;
�$� ��WT_� ��A ��0.�z�`�Ӆ�A>"{
���� �������H��n8 ���鹪I��F+
�U@�>ӿ �A�ϗ���8�W�����ԫ�>}���)(V���  ��j�A�0Βb8?M�G��o޲ ��+��� r�$q05
� `�����Yw�������� L1x�e� a�	U��t h�o��8vc#��`x' Jl������ ��0ГI��� �E˹Y� ����@�a>2� �q��&��:��?��c/��� �FN"�}�H�C����Ju��������:��%��=P�H��.����L~t`AH"}��%$v�T`^� y���z ]-3jw�e� �Sʔm�%>< g�)�^�� 9��E�4�=(���{	{"�@jFA�� ��g�.� U��P�%���[8>q� Z�	%ǡށX�Q����P� _~�+`�| ;�PG>o�gn��� 0�P�Q^����(���`�[�u 
�6�j4���C� �1�VO�~�OG���h�*s�bOE� 0� Y)�I^�� �O�x��;?�{ {s��[]z� �F���"� ,�����'
 p:�>�b�� Y�ZA�*�`Mm[j�n��i����Hĸ�`�kp�Ẋ;�*=z�+�7�G^�H.�B�;q#�۷	�x� �`X�u��+z_ #��i,������3���Zj)!�q |��I ��zi}~' �bkNc�eph�@�K�:�vV %���L�U ƽMk�5��$� Ĉ� 0���q��j{6
�֚G J)b/���>5?��^�а�H9��$��#�(CM��m�C��>� +ea�@zݷa���`E��8>�d����He0��`��h < d�;T���9V̧B>#�����P> ���xG8w����y�����+���p��@iD0�{бQ� ř��]�|��	 ��Eg�� G�(�^ڌ��tD���4���AF0B�"��E�jPڞ.�X��eW��a ���hf�+<	��ؗ�����a�Z{�Ag�����Ph��� ~�o-_��Ț�@�W�0�����d�+E(z��)�+�$���E5
�0���h΀]� �،��/��ƔnU=08�^�!��P���}� �Α�^E���@o��3a��B*�J��X"(����7�h(��硡F��"�"v�?$�hGl�:�Gn ���~��� �!��a`�ȕ�ܨ���Xs �G眞<�.$�(�O�U7���t
���V����/� X����,�	�m�D�$���$��$�T >��Vd4�(���3�A��G���d�B��� ��
�:!� �)� �-A�3�6H~���
� M�-P`0hH��E���[�Id�Ԕ��H�P�
Ag�s��b�u"�9���A��� �5�jJR E���{�p!�%dМ]�p?b>Ғ�E G|ӝ06��z0����%���	���nCx-( A�%{z˒IoT���|�m+�� q%t΅�Y����gw��E��4�Z(�W� �!a�W;� �2e�	�Õ �K�N�C� d�0��;�q\ f�I��cMi����ZSE�e�a80Pi���s� ��]9�z 8��S1�� u�@�E�
��x�)�R������ (F��e?��b�V���y ��}���C�� �����P����_p�*�H������l<�� ��]i���Q)2�j	��'�v D%����0�A�a��C���� ��g���- ��DO�����������@��� �#FM*ALvP��P�H,#/�@)�x�S0�S����9� �������H;v��
�\� ���cg=�	�/ �H����� ���%� Ÿ�~S`^T�lݫ��&�����$�Kh a��k��H$��ה�V�Ź3��A���Lj=04�D]7�<)�$UB�RFh�$: �O<y�6��$X��Q�����7�(x6���<P�� ��LHm� ݕM��ىx��,�
d(�P��Mf�`���o�'&��e� �t:���-�B�!�;�j���7����O� `����*��ֵ�Y@��� )4�*��@	�\�	6�fh?�G	%�@���4�p�	��� h�<���L2$�!��N4Hj��oi�sh�� ���Ӫ�JP���	�
���L��M�f����~g�(\I�H ����|��J	O�Ϡ3�{�E �%�_�C[g��@��x� ��	��G���N�@@�Б�3�U�1#Ӱ�H\�R�Ċ����{�:��P� .H-��&C�:ix<���w �l:nA��ဲ��7�P��ud >�:ŷ���Q5���u��8� ~X�6�i�䩑�1;�@���O�g�h�Z 94�2�	��7��]����}3u�j�1#��֠SO:��L-PA��h�P� m�M9���`:H�3|�`�X���E��"���r��F� ���=��* �s_�#����Y?�k�@�)�s��C��S>r��+k >���R�0�ۏ���*�/�S Ia�o�hy��
��\ɮ ��=� y�
��p 8A�d�i5-0�^Ў#�TI�!��+��mh�����|�b�4�1 =�K"���H�� �{*q��3�%���� >�m�d�0n�P�� �_�.5��� 8��ִ#�(3��D�� r���	<�P����pk�<6Z�0v��$�)4���I��F�3qk� \O|`xK#
	�b�gi��q�)��+С�C�&=D�y <:�M��Z�2�O� �GH6�+�48">���a��!�Ⲻ�Ёt5F$ل�`π76�|��m2�G���������w��=ZP�E9Q��G����rLl��%FT|� C�ۣqTj57��AЎ� ���"����Oj&,LP�Ā��D^M�>�j` ����O	03��+�u��Τ��}@����0�9���Ób�#��%�?$�	�70����2�%�gA4���$�iD��t���������<��?�&\ wKk�eĖ�_!�?m�����/D �7e��'��0�K�3�� �g�>��* j�K�4�i3��5+ < �V�* �a��@���N L@�hTX')�k0DA���$�� ��M�Q�:<��`Ꭸ�I�# �R>�vɬO��15�`&�|HB�1�� ��	L�0C�r�� `��(�J~����K���L�G���F�(�:�mI�d���7�-��*�"&��02�JQ��G�d �����#HIb�2D� �75�_D�	��܃־w�+��Lx��C�7��N��P���@�t���4� 1���c0�5\�����ԃ�ʹd@5 }���-Bb҇�Ļ껡���H:�I|qsbj�+�0�q��T����=��l� u�e@3�]X� Y�"S?tM`w!ց{Ũ퇄�K�<Xv  �\�n��> ]�N������6�f��z�$��&R	�0 �pD����- lvП���\��5ax?�ip �I �vPE����:�S�]b�G,��Ӧ�q+���] ���O� ޠ����S ,��%G"�� �P��NkÄ&D����� �h��@��5� g�w �T� ����1J3�2�#��X�>����`��W���q�`T��� ��u�#&���`\(���qn=���Hm��a c�(��!1EO�b�z< Y ��N��0�!�Uaj��\ ?=�!R ��X��ʜd��"�~���H�>
��}7� `��8�� M����
/� �*����K�ޔ�(�G�ڣ���j����@r� n��y�} ��+���uqj8�F�:O]����q7n�{a�͙A��!U`�@��� z�{������P�NXF�0��a隩,@ x?q-!F v+~�ҌػSp`r͡�� ,����J`?E� o!ϸ	q� p�w� ��U��e��J��b����m8�(k Co\�=LJd �-��p��1	�)������j��u?c̀_�Xs4Bkͼ� � r����\y�M���`^E��������e �0�$�su9����|���Ƒ �n�.�M� ��� QBY���� v��� �):����@����� �*����B ��>�#�S|.z�$�� �;��$e(V�Ȱ��X-6��@�>�%4s�zi ����$� ���'r��� �����Tmq�K��4nB��HG9QD�[���/���fw^<A�����D�@�|C�V-��W*�s���� @(07�±c=%	� ��'&��m eB�|�-J �H�"`���T��k ꥮ�|�%���Z�. �!ڜ��` �?i$+�c�\Y W=�"�:��f[���Y!{��F�<L� ͮɐ*�6 N�C��X ���
�+& {̉	G�p)=���/$��3���b���@�5?� �4=�M� ���̲��`�� i(%������ (�s�"�Q�� �*�8͆'�4��8HLvC rI�=uXm�FH�R���~ 1�-���n�{C,��ͻ�l�$�@�a�4����E���ݔ��%L����P�>��>�'u Mה%�W/w �}|L�Y� �9��mr���&��� �P��-�ȕ��|��aA�N��u�0Q:r� P��CW! ��2M<�����.�"p�Ba H����{�E �zO�弸Q �1���ǵK� ����*�O����v�v5L��ꀕr��w� o�dKb�v&�����g�Z��H��Ũ4�
�����G/� �\�5H ��}��� �_Pԉ � 	�zb�r�c ��ۦ��1.� ����;2s���� �� L�{0���CD9�-��j�2  a�Zb_Nڰ26��s�f� Ё��, XQal7� U���o�� ��2�A�t e�(m糫��Qc_u;�>'\�@�9�	ݙ��i�X�I&a����J����oe-(��� L� �k�* �����<� |��,�(�� }!�zj�d���Of=�I�� y���1� �i��B�[=;�F@|���#1�Cz`~�0� J5N�V:T �c�1�@<��� ������� ��U����8 rG�	`[q
<� �p���� 2e�mK��Xg"6`A#��� �.3��� �Q2[b� 9|!�j3�$:#�f�y�� xn�T�����{(! 4>Df�G����i��2 ����sv� �3�Z�HE6 �9�8t� #���i��:� �yC���8 �]O/��s 4jb�- �_^T��XO?73n ��㮇��|0���+6JsM��1����$�k ��v�WRz U�8n?\� ���1H �3��2�%>�� I���MZг�d�EyԠ��"@��x�� ���5�z� ���^�O� �a�@�� *��]g���� ؋��f&x ��^ ��K] 9aX���� �xó1 zH�!�	� ��%ג�� 6�XRi��(|�>�4�¥��]� ���
.����%��~ ����6Z ��3g���(�$� JD��۲�x�<���� 	���G��U�1����%���mn����u��`O��)���{I�?�7_8��"������gB,�A
� ����NX �RE@����9�r�k	:�����<�3� A(���6���OLK�T��N
 ����A�f; \��R٘�O�������m'p�u#� TQJ{qU��i�K����seu� ��9�BxC7 @�ğ=`�	o �H�ꍕ �<b!��w7�=� U�� ��$ o#}:6QLBO�����I��|�% �L`i�� �*��S�6`�������@���N�= �3�p2�I��E_�����J�~������� �L�(2E�\VS8�R�X�X|P �2�6��C}9�L� #_Ӥ4�fB|\�a��A�<� ��r2l���5L7�J�����K�w���ܕue��{x��]5�8�~ �(���� �����C�D��+��5������<�P�%�ƅ�)~1����%��eӷv� 3��aH�f 	! S5��x��8���2H�tX�7mྃ}� ��%Va͉B���;���!vN��ߐW��õ�$�ؘ7 Ec{�Oh �:pC���)�V~������ nd��]�8}O :=���Ʃlm��L<Y>6+ y-������W_����� ���4R�, ~�(�¸p� �������S ����,�ڙ8}�V%����]t ���&X�\G��5��_̋�-�A��:Y��r�ki6�pB]Ӣj�88@,�c%��- �_�LxSo�P�A��8�T��j�@)� �}5<��Y���Nj� eoax<ch�  *�y|"� ��K�IQfJ����x��5T�9����ߖ�0	�!��Բ��\��H�a8;˰=1��g ?���c�s� ��!l]e���V����� ���t� wySKv��E ����pj�8"P��I\ �J��� ы�d�~M:� ��O�P �Ԑ�@BJ8��pi ��*������ �A��8 S�b���] ڨO�/{Ϊ}@a[Py�,�\_��!c"T|BX 
��(ے��`��1`�z����RI0v���[�  ����f���C�S���*a�H��K �꧕Ax� LS��Yv� �e#65	 ���Vj�Z ����ny����Rk�t}��I >�|��1s ��*MQ�` ���0�z�j�!����`�� ��7���q�H�1��p� �_�j�b='s�Kx��<uU?. cA�j��d�+�r������E�u�+� &}�5�{Z������vi $6����@� �c^���.v�_O��: ͷc��"�@��OP�y� �aƛSjh� ~kU���Nu<H@Q�^�G/Wz߯S�TY78�A5C����xs
 �li�2nV���>ry��'� 	T�㌉�p �U[ǎ�@� QAFh�R� 	�S�/
%����}��5PL�=+ꀽ�� �B�KMv y�'��U�:���z�b�_|�cx�I�Ԉ��SM�F�;�2`O ��Ί��� ]�AB���-e�D�`![)�r��, J�Y~mG� 5
0�d��.҂� �=i��o ݦw6�~� f��V(��H�?�D�Q��=�� ���}s��u� ��Ч"�h� Ǌ.�lB�J�'da���c@��u �r8s�����ΰ�����V��>Te0��a$F[ (^�9�o 8m+���bW ��)���(�ɔ3LϘ��� ���I�j��c�"�_����� �Be�sP��K��{@�J+ �7��F� ��I
�i�� 6j���sF �����%y_t7~w��X ��3����_^"&` ��ӾxlQg7�B�s�H0�k@�u��S}���;pN<`ѹ�� wtu��f ��:U2���HT ZG����L
K�͛ł�����PȀD��@�@l$E$�x �'&�=>~���On���JZ\��yq������:����A�����p_&�������TzDĘ�е1��7p`��B��ód��(�
�Γ vPт�83�u6 �������l	���� �@��| �TS'���A��a0��gJ�m �.>�ʱ4YX���A��� �����H� G*��7 :j�6?�<�<���]����� ւ��N.�� 7���/� �(���ט� ����� ����,` �;�����* ���vH����2)N�9E� �f��� ���$ɓe 	/�@Э ��Ty� 馿�<� ׄn&��� ux���ɿ�� ��vٗ�% ���<��� K�d���&}��D�"^B� J��{A;�Җ�`�L��b ��1��ܲK�� P� S�L �_�:�7 JM��v�T G����Sz ϥq5�lg�<6��N��`&� �U:2�qO �IM�J��6s4iu�| �U�����	��)� h|&��
;a�Z� �-�q�"`� $�\h_��� C����� ���Tm���1֕@��W��>m �� v��\%ԣYg���5�<Dꡟ$'kd ��	�F�}�:�?�Y2d q=�"�:�:ڟ[@�&>�Y�L:����( ��5}jvƶD1IH7c`�� \���
/����̪�ۡ0}5 ͱ��E��aɚmy������ �\Jd�t >Zq o�� �s0�I/>l<����᪡���0(*�`��m�n����#=��<����۩޹��7� d-����u $Y�U
zk �<-��8˛|�/b\ ��
��E�� ִN�h�'�q=L"� >�˦� 7���q� ���O�m�� ��UG<�� 3�c�ʔ~� /�
K ��w1��d.�$m�����_8y6C� 8�
Rf @C�I��q��> ���^o� ���B�c�h TZ!�W�4
w�$^;} k��[�?M�	- n`t=,��e�1���JZ�`� ���&���3�=���:8]v�t�t�����l���r< ����A�,������b���?� �A��+���0Z/6�XF�@��< rbp�� �5��[��@o�� ]D��)TE�g��Z��>��� Ԫ�!]�*�>�( U�7� 0�s�nᔜ �-���Q� �	��W�[� ��=�츭��&l��]ǁ(wb=P����Ma3�</X@W ��PDU��F`?0n��J �Z�Px~tǳ{%/:d`/�e�@,����v� t�3��,TT�� ع���{�� ��e��g�hAR�1Qt�{F��z�[�`W��@
�B�D ��'QT8V��v/�
�{r ��x���\�^�nN��
�!b�m|F�� C*���%����H��_B �xS��(}�QQ�@�N�����f���) �ͳ���� ���iB3# R�X������ �h�8�-� +B7/��;�p T
�3�vw ��/in��V>r��B���C{R0�/ xBp�d(� ��ި��ʏX�QQf��0�B�F]" �B�8c� ����ڜyC���k@Ul(_v ��#���� ����tR�|r� p��V����x ��i\v9p7CZ��`@�.����ZkamN�T��K��  ��W!�=_J�'�G�~��w�#�а`�r����>?�> ^<���]I�7s���x1q�]H����v`�=b@����)�$�gi(UF� zNv�Fz}���: gm'�,.Խ �^�_<�� ~�?E5`e0��P�ۚ��S:�l�� щE�e��Z>�D�u�� �c^��ׇ?�s ~�K�+� ʉP�愒� �/v�1� �T����� �Q�PA��� rU,����
=����e0u �	 �ؚVC+ �02޾���� �}1mGPU\�-����.)q�@XI� �w_d#<��* �����1 �ofG�)�}��  �� D�Ŵ�`@�Bz3�����9� �?������hyk >jeޅ��� Л�>� �b��I�D�Ĺjg��*����'�Fwa&B���m6@��� ���@}��S���`� �[��e��m�X�@Z7�8��,�ҥ� /c��f@r�g���i�π�8���./l@o�f�W�6�^0C��� ���h�r� �̛�����n6��ro���E�q��c >�7l"�}��
df�1 ����c@[�3�]_�ͭS����� ����?���9�d D���
�
��2(� �VT�� Z�"Y߬��@F���%���0�CE�5D� -�ksed�Bj� �b����l �'��B�_��	po�r�1* S��:&a��
�i���tB(H,��� �^xE �b�8��"� X�{�J��g �9�w�3�X,�P�����x M}��N� ��XY�by_��c��{�3�
L�(�H �ID. &bK�Uc�� v��6��p�˩b�*�|�>� ��!����ղF y��kv$�{0o��i� (b
3���� �پj��]���ĔP.�X�G�sc$��  }.Ɣ� ��Ծ�B# $���mW�F�U�s��쾊�i�.xER� }-��#�4Uuȹ�;��t��'��a��H/�p�F&�q8 �c�4�e ���^%����&�(~H��m0χ��`'ɠ~�_�� 	J�.;�� H�G�x~�?n����Rg}��XGpd ~n5�W�}N ��jH�ugy��� �RF�h�D �Vxa:v6� d��t�U �l��J�L�2^�3�q�� 	j��/��=�x-gKW�YǍ" ��(>�� ���
&�A=iC�g�z'��a�8f:���j.�3���"�ݵ���� �Dg�'�$�{��Hȿ����]�D�G0��?�|@ ��
���� ���r�˟��Y`9O���` 뼄���~_ ���%�� >!Q�#�����_@��F0r���'}���@�VQ
b ?���"r~��� �I9��V|05���Jb�@ (������?q$���7��`0}���ɩ�� ;
�Y�dj<� ,��4iIr� �U{���e�g���!�� �Φ�N���Ȳ���H ����A���;9��,KO���G_��"����k�2Yp=���]�
��\v��n �ހb�4�kM`�x��%�x������ �G���@�0ֹX�h� +Qݯ��<�{2 i/��G'� u����$t��� �l�`n~�3k]��@�/ܡ��:�R�:9��("j�4g`ظ�͢�oi��GF+�!��;�*�i~-,Ա�s Ah�R�� ��'����&��$Td����v� �2B�0�k=�1�$9�\M��@����x ��4�ݖ J�Ᶎܩ�h��1�`\��r �N�4�8w�*�D� k��Ƽ�� ����iQnqXٍ�l3aǏ�� ��yN�_A?7���F#\з|fO�q�0u��ۗ� �w�����ҋPԯ�^ h$���B8��7�����3�G |o����LmH�����^ �~>C��	�; �䣂�ɦ���T� �ǩB:����X�)�KH�I� l�a�(��0�؀;�� 
>+qh}'��I& P�Mf19RD� ���A�����K� %k �{�����`׀[��XoA$ 9Z�d \0�y)�t��SU�� X'���]���>u��W� K:���jm�'2[J��qظ� |c3�O 瓶D+Iӥ8SuW���d��* |�`����� ���3�žG ,�M0�� ��r�F؊�?���ȉ��a����z�:�� PSn�� �X:O��� ���g��Z���04n�s�G˃: �ao���{g ��F�֝���LJ�l�T�ǰQ*� �w��� �+�r�S!��� �s0�7�j�B%��*� ��|Zi
�� ��IB�8 �P���
#�K�s� {��ln� �_���ck2�� �:ն,1��G����*�.�W���Oa�0�y �%C~�� o��#��h��ѱ��� �^D,ٸ>��\Nzy��f]U� ���z�Z�{���.�� ���x�t �;�wě' ��	�Z�� ������{�9�O �]&A
���� �vw��dp �r����%�����: ��q+P����ܭZF^ 2ÕK.��\>�i n�|_���Y�>�� � ���j}��<�
�.H+�Oip�� �X~��3�\\�) ����a'��4AD
������/ �nD�9�B ��u{Z)�� +�� �c��Xq���@�?�� ޴Ӹ Swi �K��g�7 �(��=�Y- ���+m���z�C"�n��w��V/A�V��t ��d$�h� ��cv�,�\�� Q97T�5J�Aћ����� )���5 A��E�ߧ� &�)��m >�p�8�< ���=ɱư� ��tC�� �+g�P�0y���q�;��� ���.3W� ����<�k�Z����#P '`��lA^�r���0����y�. �/�q�� �\��v� ����c&���2Ө�`���`�@� �|2��M`z�6A�ײ�h�H��]�y���O��P;�� _�rhp���9����Vz肸 ����Wi� �	K2���  1(��0ߟ�������u�J�>SR K-�.�=�}���*�s���p����X���Q ���-W� ��䨠	u��z�����4~;�"���Y�.@X-��ô��u)5� 0��h�;� ̙ߞT�u]�N.��
ъ!�@hS] ����8�t ��[̇�-G `2�<a�;�� �o]���"�@ ~���RV��Gܿ�D��K, /������ (�H�Ry� �`�/��&x���E�lp:��~ ~STa��'�������S�O@� 5��)�@({��������q���08���T��׀ACR���w�I�t� ^r)�� 
�P��t�Ŕ .�����C� ���R{ �g��åh,�� ۙk�� TX��Jiً���E�H�4\y�� ��Lj�TQ��ZXp�P&��{ �:��� ]�2�S;U+(h�� �����v ξ8V��{���]ۘ߇z�q0�:�̩	_��y�Ԥ�m��3� �� �%�V�<|�u`*�@ ŕ�a	�~/���f� ')Ȯ��υ[��04�yr�Y	p���r� �"���|_ �.akϋ	�6�qpZ^ Cx��9��	F����lh��� ����h�ud�cɣ �;� O�n
������@1��H�DD>\��vԡ�3��@���~*�����,��_������c<�D����ˎ���L׺ %WX���0$.�lX�-��� M.R� x��uȐ�Ԑ� |�s�l�k����a��[CX����� ��9T�l�
�h�a��7 !:� ����- (/%W�w�j�\�I4� �.0�7rE�UR���z����V�n�-�+8�*|
{@|�x�w lb(�tu70s�d���_ ��$��n1�M��Ip�H��,rJd(�r�	�yT���#"�(��\�Kk�  .@0ȶ +�#��t���g�hň�f�.���(6��Ts��H(�A H���8��@L\`xi�^� ��l�V�'�Z�|z� nA� Wqe�x�� ��Ш�,� �2��r��Gg:0���w~ Ĩ��R,�j
4��e��6�4�ԬX ���bv�H�w� �U�|���$�g������
�N ,�w�-	��`(}t ����ӟ��7��G8�������KS,�
Ԯ��M=���� |@�v��f^��.���wm����`�JnEY�@���r�| �����,��#(�p2��5��� �Q�����ty
)o����f �kG�!$0 ���2���ZHb,y� ة�� |> {�;��Z|U�� )l7��.�\�f��ʏ��4�k@Xqr 2�	���Kb&�mD�S�������J	X�`8 0]pW���G�M�� �y�5��gt��^�<Z� M	�2�@��
�.�� J��#c ��I����;0�lHQ�R 1w��`H����� ��=�c{�����`;�C�<$ q(]���G�;�z(+��v�P-�K�N0���Zʙ��B�)�@+�	�g ���*ir�O |_�!8趾 A��;Z�G]���c�����pI��-ў`X��ua��h0��l pU��_vI� H��e
���� 1`d�� �®g�6=�{��t @0iޥ�:u� ��dƜ�� ��2�5 ��)=���4f�ɵ��x`�L�d��������,P B-w0���G��à�.�\�PP�����e �[k�?�����L^��m� �o���l�-�R K؃}�� �7�K
e��dO`��9@G")P��h�㑀.I�'�� ��i3!�t�dq��l-�	\?�����Daz %�9Os�\U �E&t�C��_�P��h��~� ����*c �|Q[b�t��}�1�|� n�aM�d�'`����� ^ɤ�H� ��<9�� P��硬���h���6�w�=������X,�@�/�(� rY��9o� ~���up_r� ���윕��-�N3}���c<;��l�~��.��p�F��� �SG�b��y�ì��8mT xV��1�DY���,���ĸ7 �R�(a^ ��#& ��B��%J 揓1.u����6� � "���c��� ��F,-BOns1�`$+z���� ����q0 L���v����%�W�����Xc�f L�Qv@������ ��C��N/�b� ����@�{	%��܀L5l� ]�$��njIq���^�"ԩ �\��a�p��=��״��R�&"�B� E�=� / �H�@P�T� MC;���ͺ���@��'�̐_� ��?�*z� N�T�����_ ���O< ��K���� ����Ө �3o���� ��p��:��]��<[V�O�AL �ǵ�d,�1wM9s� �wB�i���V�
A�� b�8Q�` �Ǒ�[��T+�@$mR�q��u��I�@�F�f t�����^<�|r.���4�@���0]���"��Pu �v�t���w�Xo�N@߳��`�ٞ�H�1�M+q��O��co0��q�if��� k�}T��	H�4r ��U1��t+w h� 9�q��g�&PQ�� b�5������"{:���\	 O����V�� $�%d�g
� �K�}B��Q׸�ip^	�F MV|;���0Y�(�&� ʚ�[�L��E�r�O��1�.�bπ�gĂM ��^zd��\� Ƚ�`O2{+H���b�I��q���s�n����)�Q{sw1�R����X�mǫgc�A��\�5l+����.�V� �ɫv�J�2;"��1�!p� `��d>��'����$����=����;u��@�%`�,b�7�k�� �������*{ǚ��t@mN��|v Kն!�����?`!Uy�#�D1S���X<���`�ؕ�-�|Š���:��?�<
`(iӎ[W`C�F] 1>Z�	N��4�X��}�X�;�/�گآ�CW���_fq! ���"5�]���ΐ ���Bq�y���W�:�.ļEr� �0w���r�����.x�� �� ���#��t�  B�@/�i��W��-!ʡ$5 ��|�.� 7Kv����B 93�oY|��(���� {?J+B��)�0iW���m�]Y?r�_�. ��l>�SW0��9����U�P��n|z�o��7� �	%����$��W��̀0����`A�1K�6��lH�M��.���(�q��
Og0������,�K�{5a��y��Y��bf��p}"H ���K�E�c :$� ��HD�`��A& \�TV>���|yR7���� ��[�V(��=���`b��i� �qI7&X2k��F��5dGx7������� �-�eM	�W C��FN�(��7�>� ��)� �����E:�< ]zj N�	� n:+�ק/��_��u� X�z��ҽA=��`
�X��q�cPQ��Zz�V���� :*Ҋ_)L$ |-x֭�	 ��J��� q6��~���;�9�+! ](!��i�%߼^�8��
���_����p[D��� 
.	@�BO� �S=��؞	���R�K�� Rv�9���T%NJ�_�O�. V�*�L`Z��4,���P }��7̳� �a)�D�?�� $�� +��C~8���� N|�� ZV�h>w ��d�=E � ��s�- f��ByLg�pJ�����0Z;
���>��\�� 1rp�,���q@��0˵�1�� ��u�Gc����l9�x��1ɐ���~Og�P0zL��_f$�;��FR8"��w0^������b�_F��X#��hm����]���}�>u14g	���:� %q��n�AS6���#�|�U�W�l3} ��J�� �?����.��l�"q�,����Z ��͇���d�K�� ��#�e�����ԂJ2� B�>�*����NSow���~�&f�QZB*���>� ��	g �hGs�k&L�`h�$�'�Ϡ
8�ʖ�ń�xx 9|��W�BTt,0�� z7 ;'��N��:!J	�s�OW L �ʿ ˜q+@P��w�9���0�����F! ���%��
���E�Lo9'���0�X/�3p�|	*ݸ��Q@F�s֣�=��a\q? �ץ��L-Q�{�BUCW� ����7un!sl8^�2�>�8��b �{Wy�6: ~��h���� ���Ha�|p��k�u
� �Z�蚊e dF��")K�.�C��
��/���L2}&���o������N���ٝ@&3��� �#�Q�1�t:� �+	��6>5>O�;$U��� p�v��-� �c$!V�8� ��� ��`j���nM�X��萱 XiأGp� l��L�	J v�E��DK��غ6"�,b=L���qu�`�x�'R~����=�������P�(��"�P�o�p��%��� ����s��+��#�_&��9?�ŕ��
vaw��=���~G�h�c��ش\�p���CI&� ����e��v�5�?��;�|:+���g��|Ҙ�?��R�k�KTs�� ��}w�r��g�OY�6�����Q��a���@��zM�'=�h��l{pX# o7�u�8� �(���k�	X�<�wJ)�����G������>�{���MG����O �&���(\P�T0I |O��v0��җ�z�%@L� EГ0��k� [S4�]ݍ�� �<��	�V�;b�O��GL���0$��\�y 
4~��� �����:�gȯ b��\P��o�L2 �v=�J%��n��qL����|xm �u	i��L7  o�I
E=�Ԫ�%�@�Lʭ �9�T�	��(&7� �ݝ;UQO ^�5'߷����8 ��@���
��4h� ��t�ӈ9P�?�^&�� N�%V��W�a`[�'��vB�&
���"�w0�eA��1�l��h�̭�)Ȱ~ �W�ށ����8 ����& '�� �z� �fˠ(�� 5)�b���<�$�ۣ�fM�� ��Ș�c� �7�,2� ���	mx3}� �ݴ�d\�{�c]�^Ypɑ�r@g�`�⨦�H �~�ƶ��` ��擑r �܃����� �c�h���� ���S�m +��7� �e����tNî�x�H�� m�@�� r+ ,�ș�L�w ������*� �[ƻ$=��|���>��/����`�~�l3��� �Ó� �Y��� ��E�H�̓q���@r]p#��5��^�Ͷ �@�=�u0Cq��~ ��(�h=2do��;� O�#�%a;Y� ���6p�(u7��ֈQ�w}ݾ��m0���X �̷t�w��,j�H� e�qo���a;����7� ����Ҏ� n�5�+�\=� ��}7(��܇N �+P�\2��7�� ��%r���?gA��m�°`�H	�?�� 0��4:.Y� =�x>u�3 r|y�� 7��n� m��_�8�d OR��ݳ�0,�.P�E����-��D���w p����b�<�([0���Ԋs���dhX����%�A'��& "�o��! )�ÿ�{H l�ɗ-�» C(z��B]Z�� �ճS?)l"�w@<L\X ���GJ��� ��j��۵ ]�SH�B� �3�=G�� ����Pz� �(b9��q �o\�e�4� ��<EJ��w�l[ܖ���\�;���U�	���Eg�٪�#x�I����=��뮀S�� �<���3��h�w���ct� ����M�gT |����O�*�-�}����=| ��Mې��ui�0;	6䅼�V�? rm�z� �Ec��.�`��-e(u� ���ښ��[ EM��
r�wd4K�Ř	����c����� �{�� ��5�L��8���nq�C�2 ���Zc�����*�Ƞ־;)<�8�AN	���z P��t ���[+?V6 ��p%��b�B����6(x�e �gU^$�b �#����� ��	��� oLS�����ƪ� �>p���:��	S ���= ߚ��`��!�e@-�\��� jw��(L3 ���a���%d� ��c�ۓ �2@�.��;������X7 ja�v�Y3 ֲ1�sHC&��hr�� �'jؾ�mq� 02$�x^uqw n����>H� ö��|�BU�<��ߠ�I� �d]��/A �����G� T�q�EC� ��z��Y� \���±��+
�ǿ7娘\p4� )Q��� ���M�t�G��Na��k��O��� ��pz[�U�`�@�(�� D�Ήm ��d��RY9��P�"2�y�� �:���C��&�L�	u����
�Z �<�wQ֊���|*�.�ϴ܆A ���2�,F'sNn���/gi�>ȝ �H\�j� �����7� x'��f1o� �W�%���h;wG�v;�<QV�j4o�(w\�<�C�� �3 ��D��lA� a�K��W Q"�?FH�t�l8fc�]7��&��#)\�z �}���O�r ��P���7�ql_p�d���g �:�P�( ��%;QÉ �y��$�r�.>|M �b=Nj �y�Y�J �u˩�� �G�P6��R���Ov`k֛ 3b��ƃP �ܘ��ʩ}�$3m܂�q�\�� �5��C�ے ���/��
V5s ���W.~ Ff;y��}s �W��� 8k72#� Eb��m�& q��?f� ��2r��>(RǠ��l�&��J����-� U2��Y��� gz6!��J���	����+��QI��� ƙw2�=�� �+R"d��*9���� T�zV���b�O<+�g�ۘ�>�c� ���ly�;^��(�T��D�� ��L�_7��Y��z3D�gX�  ����J3�:c����K9� �OjE<� H�ꮨh�� �'��*���ӳ�Û���J�!>�� ���1n�Z"_x�͚�[� ���|8I5g �]�T�ف	}�3C���5�+� ���kg_� �M��#Fa e�D໷���j0� a�Hrɴ|�<�Z�Ƙv=�\ ,Aw��&���ǈ�N�v(�6 ��|�Ǟ�� o�"tV4$?T�x
s�h �cA�$K� �y���� xS�RK&�@���Al����0(���������`����!{�U���T��.p�H_a�ĐL����{ʌ &M�087� ���{�IZ�h�g�`"��+� �T��佊 ����:X^� kG.��>J���� ��1? ���}X6� ���#�E|����@�� 6:�wŁa$H�z ��)�o������%	��]5�w ��sX�h¨gR�z@�`^v֐��w���YrTN�� �R9�5� �=Т�w� T<S��ԟ?s$W�mޡ/3��Yn�'� �zf���~� ��
7�	���ؔ m����ױ ���ɿR�ۤO��o� @	z� ](�Z�^6� ��9|\1D�,��2aQ��%[R1Ů �G\�c���XQcc (�=��F�9 ���:�X��&Y�t �7xL� �I�pe���2� ۛӞi�� ��J9}a� Y�e�@]#> �l�\�;�n��2M ˝���� �;�nXb� j��Q��� *z��W� ����2{�|��m��;�,% fc�BMZ�. ���A�� ��r��`W���
�c��.��K�����HL�y ��pk�De �u�&�s)�����Z�{a�Ȋ �]���$^51 $��`�% �P�a����������`l �K�1*�D Г�b�'{��� _	�M�i�(� �Z��p��E���
K���Qh군�i��@��t���gp��v{�mHʇ��-���E ���CV`8� �Ǧ?l�� �p�=� ��
;�^ ��MyZ̗�L3 ��P����ׯ�����D� Ƭ�9{�	�Xn��� �\��
��� �����-�Q �>ڟW�x��+ A�6?�_���(���i� �Z�p��^�`�<��" �~�����*.S=����ԀfG� ^}����4�� /�K:A>z�l�%7�	��]��|X�M07��\�@��X�S wgH�����+c8����� ��$�o-� <��@P��� �j�i⥝ ��_{b�� ?/�K��� ��`��-BI{f ��}�0 �Й�^ܥ| H��?ɖq��_cP( i!�d�$S���F|] �Kê@. [��*����P<�h�H9UC�_D |�R�]B{s� �q��y����X���fF�u�p����K�b���sf��U�wP
�0:�� ['������6~����B�� 1�r8��6��˳�°�D4oҾ��<��C�qB4�����?O/(ѹ�������q��L�u`\�5�ky �{_�7�z�t��,�T@���
�m� P����ќ@#W�n�IK��b��X��M����<(�/T�o� [f2�#;�� 
�'DB&�m<�z�u� ������ t�x�"�R�=O� ���©J8 �\7�y$Tf��"���9 셸��� �? (�I"�O�� ak+����\��:>����	�i�H�H=1��(�8�B� ϯ��Ga�� Kqf�C*�F���O��TQ�e�� �����x����B����{f���W_��/�	ߏ�C����`�������'k��� �_2������ �a4):� ��,��tF��x]�ƻd�����-"��9����v@�*���7����� ���c�>���0�[ ���H.���{dÎ����2��� ��`����M v�!�ޖ-�c0{� ��=e�J.��!PO/� !�Tύǉ�VZ@`��`���0�'u\�Om�H6���h5�P��� 'T.H8��[S/ʥB2��(�� ^�P"aI���}�K�H"��w�(
<:��؂ȟ�Ɩ�-ױ�P
�чƴXo|/E�(�~)���`_�3��Qh�<������[A�$#��2m�yb�&ca�@����
���Y�p�<�r�0�b�+�鬀'�ڐ�-���JL3G)�h�	�(秡�\@�I��H�(,�4.�g�(�y	�z�&By�\�v	�~��&p�t���p�L�X�@c��Ċ�>``�[�Ic)tb�l�3��Hh�x�7
��e�H;�(|*
�o�����,Г$0�$�W��`%"nj`�D -��5��LWdm
tL�D�=�S�G d�������<�9K�oJ�@��1}wx��L�m)�$��fh|>
bT�uԒ��g�����LhS`�Ww��N�()H/-�(��uZ�	�ҁ�k��� �կ�e2O��<��������8��� (D��:�pge�@���ں������;A��G�8�=z y�X� ��ӧ�`Jf��x&*<@RI�e ��Ӈ�Y���:�Qa�@�g$i	�,ǆj��a�� Gp#J�v�F�	�#/���'��;��G�!�XPey�@��Q����P��l=�w ��N	��'s���_J��:<���V����;�u ���x�� ��ZV�~y�)2:�bLG��m�P��dJ�)�_�`{<�8`�0���/)Ι,���{��д�;Z1.��&@�R�D�X�(��B�k������I�}d��\͝ |�_f�.r��e=^(�Mi���mD<f?7`�)Vx�����/��_�t�h[�x@ԉ��I�Đ\"�OYg�7n]ER��Y +6n=� ��?(߽�ay�Fv��J�@u��_(��1q�0������D�~.�`�=F�m�wuy@��H���	��% �|�ǚ$f*�{[��cn�g��<tЄ-�z1 h~�n�ƈ{V r?[�:����ɇ8��HB,��y��.7`�����DߓX �>ty0H@{Z����e��_�8`y$0
dpHk~y?2��}(�ذ�O!]J��J�$;���=��*��H�T��0v0 
Z��͘��K��G��N�D( ��j�>X4x�y�e?��C���������$��0n8�
|���9��	U$�✼�x9� 4��
�]�	U�?�4,�F�����@�@��?��};��h$go4�"�H��!a���h� �}�<m���o*�3�@�B|� �Y_���� �1�}(���?�YM�(ѱ�(���^�:P`��]����8_b��c @鐃Q�(� ��[���Lu3?���`1�����y�)? � �p�|����
�~�)@-��/`h���1t��y�`|�Bd3�	�aZ(`�h /�A�>t�SiP�Ō~��jB�?���!pA�� �p|�������3O�(\����+�)D@�׎��DE�y�𺸄��0h�r�����L�`��"��/���P�I��ϴ�(�;*gZ0 ?E.@,����	���k!`��ьLH�
V��z��M��(��e���(�r��%^K�`�0?׹�0����u��`v�<�dL@|�<ہ��J�0t�J�2.N6�i0��x_�(`�(�fe�p`HÖMg�I���{�8�Dj'l܂�(,��a�~�J��
.S���| ����(���q,���@����2<�V���� L\��������l�1a�
�<��>𖼐41m��`0P�	6�� d�9M�)膰H#P�0�P�-׆��`���㨠ܻ�K�P����a^��z`L��@��&�
h�,Q��+�ڄ0��86�t��\o� ���A��4@�VK~�@���	z
I6D���㦲@�`����u۽�A�� (P���$1��#�t�Ë D��� �c�hO���q�@l�ܨ��܌���~`���GK[:Y�����\�A���1�K4q	�Z%L� �^�A�:@z����=��P��.���~(�(F� C�}���K���dSϘ(����Leܪ�����$��8��c8h�'��(C����tz}K��Ih�	?�����1���9�g�`���� |S�MW 0��G�ՙ�`��4<IZ��� ָ�:�@p`�(���J���( #� T;Y�p�{S$�4<�H^R���5�퐨|��8d�dM�+$+D� Z>�,x�N�X���E©�3��ބ��E*� ���O��䚠M F2�^�f퀗�$~���H{�����2��πH?y}�V�D��B��X����䅘 %�:����Q��"@���7^��:�	 ��q�~�옞aP� ��A>j@~ �1<H��@CI���~TK��xÚ�4 U�'�c(! 3&�-��:ҭ �;(�Qv|8��$�1ԇ�b'��Srv�%�8�q��0�� ���!p�H>X��qI��(^�LC*������~j|���F �"ͱ&��`U� �)!�e	�����(����v��1&5�f���a�������XB<�LtZ ��G><z�'uq�c� (�OS�>\P{��ck���� #� m4�>|���^2�0H�� �F>�=&��0,�Y=�E�мc^��+(���<� �_s����2)@fPB|4�إ�DX���O%�,SE��0�e�̪ap`���.({��(����]г��-ŀ\����0Tۦr �?|wQB�(�i%(�����3Ba`'JXv�ؕY��r$u�XQ��0{@81�+�$���&pv�0�8ހf-��ˊ�dyj�2Ӕ� ��]�k�� 
#T8'�MI�!�G��2Y�$.V � G�k7�h� &���� Մ�T�0�R��p� &h��M� �D5�ޅ���\0�q�hY ����u�\ ���e�� '�gJ?��/bܰS
E �I�h�*��a��=�M���� �׌��x� +�?�i�� zՌ�{w�x��1��JA �)��ǵ�ne3���x�	-jp2 Tu�p���q�P����g� Q��ep�l %��+����J�� �9V�n�$�b0@�>��! ��Ko<D��%�����# �$	���� :{�Z�� `L�9��f �h��W>1q��7VT����M�Js� ��q�r.
 H��NM�|P�`o͕� d�r�*v� �&:�b������\��3K�m U�}���� �k2�tl|���n�"�a� R��J�̀�?�<����V��:=O &��Ic m�b�Y�� E݉���x �,`��.�1~�`c0i�grbJ��S���3���GQK��,� �s���+�<���j�P��u��]T�� �!J���#w� 7���� �d�[4� �p@��玠ȷ|jRu��>`�  �^��� U�ӕ�W ��*xr���z��)/`���Rl�H1��h�r�e�i7��#8/���� XuIC���x��/��.�� qLD�������1# 	��� '7ẗ,-� �&0���ňL�̐I �qMo��/���5��|���F�݈�U��ј�c�n�l� �:�,�-+�G��)ް��h(-6X����.�?v�s/ D���u= "
^����`�W����B4 ��<vjc%A�V� �Q:W� ��gB�4�� V}�1b'#��sM".�� �h�_��� �N/ђ׼g�$�v��ç>��0�SM����T�\�%�����N C��cS'O�@�@��	 Wt�x�s� ��
i�1I ��%��E ���"��r�03a۩����^	�*cz��4�$G	`f������H�� Bɸ:3�<����Y�̛hP爥x��E�BI�������P�d����k�@��� D�U$n=�S ��3��ah B��]���S`�����q է��5�A#��F��<
"@�3�� ۠�Ն Q$U����;� ���73�8G_��5R� E~�F���b�'�c �i�. �������>�q*�X ��H-B��@!]@�a ��y2��)����9pi�>�.`0!��� ��(�������Lum�՝�  �\n_��� 庠7-�=)瓈%��6��D��B����&��5 �VF�=9� �"3e�ġ�� ��V	(9����qqtL`7��Yp�&|��A��PG c��Q'�Y^��0�� m ���&F��Bv+ �\�cޟ߅-���BP�R =��5�6�\��@�J�j�� �e�)D� F飮^rM�io��W_�
�L ��f����4��`z��J#����Hp� �S.�� Wv۾"����7����]*r�yZ��Y��i�M ,��"�W�j�P��|b��N <Ɛ�+�X͆�. ���^ xI:�\�_ʎ6�;fw�i.�: ���y?G�۳�Ծ��fV��[��;��ot� <�`JEl�P
b� ���e��T��& �%��������;B`^����[�|g?�	��A��s�/)<@z��S��?ό��A���$F�a�Іc��������cS@(7�:��� nI�{��!Mr����� ��Y�P��W *'dg�>@ ,���6s\�x.ϸhT��c��/D����n�Vs���ƲD$�@�1y�00@�`"#=3�K� ܫj����I�PF ������a�X��/S�@�k�t� 9Ԇ@�Ǐ!J�X4ڀ�
��& `��mq@�O�J |�W�� �|��ῐ��>�X��$��\���^�@�-WO C,(D�� uB�`q.#� @�4�T�3p�C5�ك����(@�O|t� �E����g�@+q�` �ed ~�kuhR��+� )�W�}�Z �-��J��y�&��M� �H'i���Gl���=��bj�`�U�Ǳ(� ��n��y�� ���L�{�|�5o�@*�nۖ� �_�
� @���2A}�?��ۓѨ��D�|� ���b�_���5ۦ��B��8S�}�������wّ��;��K$�w@��J`��
w*���`L���a���� ���� ����v���y�%� ߽�K���V�zO:���P�� З'ᡴ���X�� �7D�py|�!�Ya�ׇ� y�
��@Ps�uL�v�K @"s.Q:�À|�WF�`��Ov,x���NH�@͒���g��ダx�J�ڷ +�O���� ����?x�73�8!�} ��Eݻ)�i ��@�8 <���z�g�>c��ǐ'I� l]���C� &���?o�V�5��'8���9��3� R�R��V�2��^���P4�}_�Ӻ��@��
�S �|� l����!� ��<���z� .�Uf��Y�� ;��3H��P�����ЋnGX�
���
(JZ�]҂D�(6{�9$���c�:�J�ǵ|��#��@��`���������GQ�ބJ Prw2�wB����
�o��*$!��@�_��# I�r� 5��ll@n).`��_�E�`�|�rVv@`@+=�FW���o)�@���E���@sQ*�/�$���T$��@p/W��"��!�`]���[@)ƀ���G�� Q2O�۪]���&b� S@].���`����@�U"�`����� F���>�� V�qщ�: J4"�A��Q�9���
�n@���=�� �o�����ʈQ��-/  Ox� ���g% ���&O�����8�<�n0�0�R@[�.�B��x �]p-4��`�P`���U1�� )�� �Q��me&s� �×.��R n���=U(�{���;��ǟ���w��ŭ�p3�Y���������h�@���>���b ����v� ���d!>�V��(u�+H�^�#��@h�F� 5��g��,w��kӇU�n7ܼ���W�s�H�g dD\�X>b  �����S; �at!C of̤g
������W!���G} ���0:cam$�\��᩹�
���Bj&r�PI�@N/�9t;�oi��Z��Ӥ�H
�0���] u�4[��ؤB���� �O�D*h����Д�T�f,�Jmƭ��>@����P*����aP�K{����F��,f4˿1��P/�� k� �j���n�0t�/�����v��ɴ+-&x֦��< ��w=vh�����%�+]��,F�I񀐁-{��pE  d�)� ���8��/ �<�� )p��r� 
�Wy�h�~��& �$�S�<���%k�VZ �{��<��V!li��d$$W`�HP3t % �d���"U�0�$E�H�45[XG�=`PS9��TjL��aCI��穗�+�BJy�<�� �/�L��P 2~�u���5 ���@��M4 ����L�N|���O���h�e�9qY���=>�4� "�H�3 �ԃ�]�:�̅U��̀gr�3 �W`(��N��|*9(�H���(1ݰ�8�%��u��1��,��0o���f"�3�OU1>jZ�x��"{�0���հ$B`�`$�V��:�H�瀰&L�0�.��(�[�fu�X� Q*���O�y���Hڏ�\Lp]�ۢ��d��-�:�� }��o�'������w������-o #��:@5� ��݋FnM�*��<ܘ(�DWa�ͼ�p/��W��s��e���:�i
M��<��a	�!�i�@���x$d�<��%�?W��&�m��:ۊ1��\��%��� ��+,�Y�耙�1L�@��0}�P��~
����`@GK�����0p�@���g�#7�k`�_-����<�ǘ����H��by��Bt<u4��P0Ұ�.�ː�
�o�WX@ywQf���CnX�(A$��p!D�x��g�X��)�ޔ��j�eY^���67�1(��8��T솑B�k�蕤�b1���b�1]L�T�lHS��0�`@?������`��R!�{�'x�0E03`���:��S�4�Bt��8�B��5!�Ϥ"�0��L�D��L���B]���e0 <8쳆*P
xg:���p�B����(n"����䖴*'���`I�P���r�P/�:�0p;@���D�nlTAs�T�̚�>�+��
I�0�����(p�)����Ė���3ؗ�a�T#�&�����[x�����i��8�mԷFd,���nB\� �]X����� �Ǿ���Z�˔�G$:~�IeS�j������0�di�����.�a ��X`(�@�F��� <!?*n���#��p0Hm�XT��?~����%M����B҂R�� 􅫁�q�2P�`��Ml&�6P�	D��� ��� �8�M1��৭�� r�]���Ű �1�,<i�l0qE��xk ����@�a St9*�1#+`T9)�ϐ�7	f@>˼�R(�uehԮ �s��8\��AP>�3Ђp� GZ���/a�P�Ӌ���?my&2� �9�g�oO�(8 ���)hiG��T ����C�
�;	c�?.�=l� ���Yb4(>[o�F0D���A�t���0�V�z����0��u�� Q��+`B���[?�R�	�w� LefUNP�Z �m�c�!?�G#�9/ⸯ ð�]� ռ���I� �?�0�H�O ;5	��q��di  .�OK�h�-_��(G�:4&��%A�= Y!W
�*h�+�����L\�)(�q�
:��I��c�fd�B` �j�HX@Ǥũ-%送�QZ�)~AT@,9ձ5
�|Ħ�}��� AΔ�6�T ���������`y���[L5`=G��@q�� h���s� ��%+�}�M�3*5Zd�����
�xm�E�̖��YH��O��$P� �
�ͦ���k	�x��T�$b �B�C��>�P�H|@�{�:�r�H9� ��*q$���k0I�U��D�aw�1��-vN&U���bl������L:�&��G��*�<�o-	,��
$)���G�j�7�,	q:�t��"����H�!x0��ӷ����߆�4J�4��Ý`���qݍi 8���	Q��0�} �*B��%� "��j���}��v@X]O khW����Ò��"�
��p� s�I9,��@PX�������A`���`p���a�j%��������B�,��hļ�=#(�/�Rx��k�!���=�w�$�Q���Q̈䛋���Utu�0��@���E5@ɰ ��@Ai8~���C�V�mE�P��rPʇ�W��-�e�����0P̙ $��5j���&۷h �띉K�@����8 d��r�-� pDy��1&(��=Fd���+f�R� B�E� ��qO)D�2Z��pȵ,08n����BR�$�KDƍ3"`h^r�7p���F�s�пi^���fpr~� ���k> sj䗿�e�T���0�tp�?��4%��F@2cs���6H��t���� �Nv�\���$l*$�j�>*����&r;�������_��p�Ȁ�I i#�ˀ���NZ!_�;��j@�|{fa�P�{~�@�0qYW�]A�:b� �O�� iP 7��R�������B@�E�c3�\o���_&y00E�@�� W����;7���Q ��6<!�-:0g~���@��� �N���8bA�cr�n8����S�"�`|��-c�� �8J�;b� \xq��V�T�W�!�4j�T�o�0�� �(�6�UD"yn�����5��x� �H1<`3Ґ�� 0��� =(�w�T�d ��Znܟ����#�}�W�̌��+$�����Tg ��o#[�_ ���V}����Bk��C���V�E@��ם yżղ�G ~K�2�Y����� ������� ��MÒIv|w[��A���4�3���O��7א���o�
1��{xPQ� �HO����_ ��n�]���� (+jF�c1�� �>C�J�^� ���fv��U�QX���
&b '��Y������mo��� �!��"� ��[N0 �?ߗ�+��Fsj�����a3�� �(`ߪ1�R Ң�H���$��.֧�UgP�� �w��p���`R!59�`*p����90�;����"��W� �-�5�/�vH��p��Ю\ ��=�g�> b�*�4 �����P"Ce��*:ه�k!�h�q �(���CͰ��/���A�̜����]���y�� e3Bb6�xz �.�)�� C�{�qW!��襀i$T���Q����-1�� U��i}�O ������y�̰�_q� ;��i!�� �f��J�c��������*>����ast������(��� '��V繞�`�a^�bҐ��ڣ~�9���(w�L� p=-���g {f�3(���� �UP�4`刭3����ab�� ��o	��	��(u���I՞�3 �<wf�0�7��Dg�H��l���f�;k��(��� ��v�6�E �-�',;��ݺ��à�8��?����aG���� ����f,�l`h��
�b<��(�4 ���H8T��x�*z�(�1�.�Ҡ�:���h�A`����c9:��X<nW��d;%o����H���.� E��O2�0VbDڇ(AFZ����NC��q����=xU7������'�������p`D�'G�3��6�C� mY���1��I�gz��۔�>�LP�*�� 0�t�W����} u�4��Zg�320@���r!��ut�( �c[2��>�
Eۚ���FW�K����_� )Y#Ц�$ƀ:�Ȕ(f|8��(d�e�/����Q������\hT�p ��H��E)��zvc�ȟ��*^��6z�a`�P�� >���{_��pc�H�� �,x���l\�� /����K�H~ {� �?g�J(�s���9���� $�����>�� ���	e����pĝ�~�&`�3"@/*�� ����,	<İ� �0У{� �~�Ȭ�U]�%4R� t�7% ԋ���@� |�¸��, 6lb��$�^ɕO���nEP�|�"��q[D�A!��op:�ބ�N �I<Va��ud��`{��0�oƻ��p�W� Nv�J(� ����~ i����kL��GQ��8 ��πL!������'�йE� #�9L���7(��	,3���<
�~ ���y܄��)�J�)� �9�*d�7 v5�n^W ��,0���Uu����L���������CeUP@qw�r <3���ve�7[�`�C���g��d��� ��7�zE����5�d7\M���, &�f�3�yc �n�RX�J� !-%	#]h0ـ����.� ���{nV�Gq� `���R@`��=�� Jsga� [��o�xB_4C��،me ����_Xd�v�v+���@r��]�� h*�t �b���>���0�] ��(@R� �9���3 �;�C�- �!��8 e�m��Ctb Oɨ���9�I�����/2 �����k��]�׀y��, `ͬ趌�F#�L���� p��t�s�		u�K`7#�|���z����|����1�]"� �R��x�H٭�kh��l=uL ����,� �/�\�ϋ �H7˻�:H�� ,�%�8uP�Bh TWA,�* Z�R<�� >��l��2E�U�)�׹ P�SB�0�m:l���{y ��2�U3�� ��)����oڿK�#O87 Mf������Qpy�����y �U/���IȘ�>�� �G���Y ͍�!Bf#� pL��-s������P �>�K.<��� �D��5�{t�� �)̓�\V ��T���42�lNIg� �s�[�L�V=#a����%�}c= ����k&m�:�9^��� -3V+��}\ �rp]F��=w��mz�H� ��<�B�r� D�ߊ�� y�'e���8	d w�|�cqX����R ��'��D���[,���`��� P�a\:��8� ��˘5R(1�OB�հ�8۰� 'ٷC�� j�6,@�N2�����M<{*`�5:�� ��/��A� <���yU[j�N�5d�c �-J��R�z9�� �N7fѨ w���D��  ���_s����L�r��[0 �}T��@c�(A�?�W�Vy� �H�K�� �'ہ�Wn� ��D��,:����sGŋ�4y?�uT� �1�r\X O$����'�ȗy�Iw��r2� �]�Sn/yw�"�1���e� Ĝ͇���������������ȯV SP�E�+����AfU��~�䕡:� c�_R��/� �������� o��z2S�V�u�� ���r��� �x1�T�6 �&���ۧ�La2v��m(�׍�{\ �#���-�5=�W����ҠRo 3	�S"L6\�Z���_� [�P��,�{ ���|im�0�/E� օt%b���]>�a�(p��c� �J�#�F��k�$
�@:�� y��rWڜHP��� Ϯ�k/���(��p? �]����1 @�r<���u�=4`�_e'�$-. �D?��\ ����7/ 8߽N)��¿X$� �Cw�A��Z������@�B"�q 5��S�� G0Fϲ�EI���&�0o� p��S��t]?��}8`�wĪ�� ���C!>��0Ҩ�z�.2X #�ޖ���� U�Cɱ��v ��ߑ'P���)��G�]�u��>0��!fy�9NIW�� �\>B�z$g �8D�*��l0ΕA>-�������@�P;���(���*��ʵ�l!��IԠ�=�q!"l`N��,�:�x��^EJAŀб� ne�� �aG�A���K`SV=��ǉ�tP� �avRS�X ������� w��#��|��`z 6�i8MH ���o�۞7f}��°{� /���1�� �~�7xW �uM1A�Qn���~}] �9��V Y(��BՒk����3�� K��*�fv�\ew����@p8;-�1 L�A�À8� �"ON� ��EXG	f:.�=A �����/)�� B���	�X� w,\k슰ҕ'��6a�# �Xt"	��w�zY�&2�`�sLZ�8��Q]:0���L���@��& ח�_dk�� 7��/X�+P pCQ�ֵ� ���}��&M��w�|���R �v�Q��Kh �ǜ�;�)� �⓯����Xvh>�83p��G�asNQ(�n���!7�>gY]e� �޴�0m� ��#���LnX �1�+������C׃Fl9^q �[���? ���bں�� �!Vި� ��t8���#<�a|������jd�R(��ELO �S�"�4����y��$��p��Q ��i�̆� d��>%;!� ��A�?�L8 b(�-%q�<�p:|��v 9^e#c}.�s���C���@<H���������f��� �IX���4���ZO` ��ʻ���L��߀ s2Nk*-` ��
jt�#Y 饬B�Qr�);0X@c:���$�L�_�P}��D��I7 Oy��8�Y ��?��Ft:/ <^(� p,��Ӊ�u9�e �|����R�:x�u��#�C �^�B��> ����S�[ u����5/��� YV�r%��J>T� ��  �0.q�����Z'�����>��A@۾b�&^ �g�2�n G-�·b� �z���=Џ�8�@� �v�{ �qm|K�9f�E�˭ բ��#� ׺�1��P2&���4�X��]�+����ɉU��78�
 r�������p5J��Ė� �7�<:��H��}�;���e7�I� �C5�� 
Ժ~�x M�R�=�������+ ��>deb��)$��J�h�X �3������ $��4��.;P0�fȳ�� 3��?�{N� ��c���)b�áy��+�5��-��Y��$z� �/S�W���Շ���j P�0͎�UI�� ���ؑ� ������]�Z�� OJ�&!�S� �r$p�F y:6<�U� J{wX#^\��r3$Pu��J4�n� m��B�S��1dG��� �<�[l�� �R�DX� J5���#P�PE�H��Q[`�W��Z�vn���� F\}O�XNI�#0k2Q^�W��pB6��9�+ �{��u���'�m ٷ.-����<䔀�Xz*T u�)�YIM<C� ���Ko;:~U j�}W�ҁ�t�{ �� Z]��W���K�|��K�"� ^��V��� �,/�A��s;�R ���|l[QtJ��ף�M�D 0,"��h� ;$��B�� #�&]���� �����
+[ T/�g�Q��X ^��\CK� J�8՗��� ���N@����V �q0�J��� �^����' �>��ԁl��`�� ��	1�vR_ �4�#��z  ͊߮�3 uL��lI�<A�BJ�i�f,|DO 1}��N�@��F-���YR�@�X��h �V�6�B.0o�� �<�$� ��V�ɬX��2��[�?J� /�zLح�� ��	�!?q":�(�רȯ�<4x��a	�-� �L1e�62 ����lM�`��D
����%eI�x�����v ��ݲ���9�� ^�4nQ� yY�!�s��; �$Ee���<� Rz�� {��qA�� D���e�� f���`���vLݴ=���� �'��ۑ:I$?�2 tM�K�� ���j~��p` lW:_p�i�CI��%@:�7�@(�az� ��\#,�w+�_4 .����H t�f�	�> �14�LM� (_�?��}p !�|���� �����m}32'~����� ��A�u�o� �T�Sp� ���6�g�	�F�Q�C�El�[� ��.)�1�N�ƞg _�C&<�� �U���fL�^]Q��، ��� qw�"�h� �Ω�]	�g �%B#}~'�X��bQD�����+" u�x>�4X �M���̖�0�^�>F��YO�1� L�Q��� �2��bU��OƗ̢��s�!���ޜ����U(�]Z ��#/��_7~`�0O�r�p�(P���@�ɤS$�)tb����q��xK �W�VO����?\ ��7����K`i<����}J� ��X��OI`j�H�htL ɷ����n���T�޺�� ��V����ت~����WL��R ��U#�C �(e�EI%P����B�X2R�i��R ������Ԗ}W��r�.p�:���hӊC3��Ia>�+���Oi~� ��e�E&qQ2� �詑�"��?����N�,�@�u����3"�8t�Xt�Hֻ��Hrxh��� ����� �B?�- `����y �\�Z�L� ]޲F��a ���4d� ۶��3e�y z�fCc@� ���'�����A ����dj�qr�\�x�]�m�p� ��\�C%�� �{9�I�a: .���\"� Ǹ����(�}���' ��v0<����z@ �5�dC#� �+���� �$߈�8n�:B⁶�oz�`�P �!�~�r �<} ��]* �۳=��L� �!p�Uګ ��9�ӟ 8�e7�<$* �u������=�}��8F�$��� $B],� ������:���!f�<�}9 	���w� O��?�~}7 Y�p�"@s_ +=]6)�d�a~p�_�=-�,F�Q��~ �3E[��R  ��סWL��0(}�%��XI��� �Ha�/�� ����NP�}!�o�a��ܷ<�k�(�Q�-3�� ��{���g��F����N �	����������7az?�؞%�ꡪ���neFخ6׻K�����p]=>b��N��,�WUz��4yR��E��w� u������Zw�^O�bɣ�.!��ޛ��h&�j? �ۘn� ��d��QB� �\U���# !�(G��� �=r7�4� ����aR�#l}�'����� _�LcV`b��M ���i'+�� Z:��t��|�01m���j��Y�����wu S���7�{� h���֚� e	��&]7Z%E���8�ۂ 3��6}�] ��^���C���@�`b�u4�<h�Ҙ�ӌ ]u�=�/��%����w	�(�  nڰ,r� }:R�8mE B]�4����+�q����� $X�dWѓ|z���(� 1�e枴�s�� o� 6�^g��i3����Q1g̙f�_lӔ�Ѧ�M�E� �f(��
|A<�^���it�C� �m"�ѭS�P�6�#�\j��O< yhp�z�m�zl ���͆9��=�G3�'�p,]	�H5� ����; ~R>���y��1 �a�N��!  M���]l �
��:6�N'Px����a �7ʂ�z�<cr{`f8�o���9�� �>�b� ��u!��)�����`l�:�E���T��� dm#9���;<����˥��� ��פ���t���z|�cӿ �d��i��@s;�${����o��Ҹ�`�� �^IK�Fq�<%��e�L��mҖ/�`Z�A ��,h�
&T�s>#dþA�)͞�E��6�-� ஐ:����Ϭ�L�nA�c����� ��@7��2���*Mܓ 56,J� ���l��AyΊ�`�Pǡ� +��`r�� )�"v�yR�q�1 ƹ����� �ҦB�K�:^a�I�(�{>�Q�غ.������a�;kJ��p[y��N 1;���G e�ah C\���ݝ�X�Z&f*���$NA ��װH��)I�����[ 7k(y�}姐�9��z�����#� c�{n` ���;� g�����x���x��z�Ě l3X�A5� �)�"�Z�<�:�F@�JHg����? ��|  	�>��l �Nt�R�a�e�CE�@�Q߫w��	�*ΎI`�Q�!� J�\䞃��@y��� ?6��(.�/\F��= 2��h�Xq ��<^��} �,;�%vd��?�u ����p��A����`�@� �J�bB� 7v^-VY`�S}G E����]�= ����>�� z����GQ}8��v,f�����C�� ���+x�'�#ň���9 c�|1�&�{� 3��.CpΑWks@�M�}� z����	��� �h?j�/�#k�%�����
<�ﳍ1 �����Ʉ0� ��˓�VI�q үݪt�x38�Ǐ�<��:��]��0 48�eb��daF-����+,�� aE$K�֟pq3���ّ�@p` ���	CH סo�yOR�q= ���/hd��q+��U@0S�����d7Ō�ê�j�,9*��\g xb��28 �(�u7�.<�� E5���g��ڹѽq���8� W�-6�L����+�� :�?䯁 QΔn��T� �ЫӚA �=�*��� m�tj�CL GV���0z ���dvmNPҌ� �� ������ ��cZ��Х`x�n�� �h�W>5aP���P����q41e��3�L"�� F�D��( )ʴ��9���Kd��L-�`�XVG�\{ܯ�|��n�^^P@G�Z�!��� ��%���_  ����� t�y׼�̤ ð�I�RxO L���h@j �{�!V��R�3��6  ��K��;� Ah�I"�� V={\-��&�˯(�����X��p.?� F��n�Lm�� � ��
:�wa$�L� �<�1? ��nz��K Tt��䭩��;;�|�p?��9о�� +�W� -�l�%���A�� =q�[�6D�t �W����>Xa���"�;R�� �!Q{�- �	΂�~ 6�w�"<vbY@�
�?� |�����Vhi*�HE�0�� �<�;�50 �� $�<�?��Y�i�Gu� V0{*1���C����Y��3�r�����z1��{������b�)dl z�B����G=��X�Q5�[�7� O���R�Y>�C �,��`_��� ��Ի|��L /�y�3ߐ t&ɳ���� ��8��d�� |X����&� b�q�w�'�QXf�+�,v��D�-�Ya�|� ��l���� d��_�� h��t(� �����ۻ� $4�O;7�� �K���B�� \������ o��V;= ��w���UK G�o% ��Q�0 �V~��H ;�/9ĝ> j�4A{�F�&�7�Nk�`x<�3	��
dm r2�6�J-(�	p^̑wZ����h B~�z�= �����| i%W��7� ��.q�Z�~� _���|��o&��� G]59Z�@k �P��B $�J�в��6y"��_ l#C}Y�k E^%4DT��,L!jo�$�<d\��&�������$~h M��P;J����H�`���}��j5 @v��^.I r�c3+U�� ;n���v�Q�
��^379���   �[l��� I돼3�� `�s��Gy$X�d �m��� H���}Z�dY�O�i�I��
�"�� ȶ��u��E�z�4�)�<C�&�Vج#	7���>��������pM�� �^���'��qg@$֍,S D|kҵ�>���[��r*?�KS�ǣ��7�r y�[g�X�&/�T9�O�r��(�Gp�m�%�3`$�ۘ��M��:�(\ai� ݂�	w J~���F�, ��ŐR�L�⾱C�@���� �t!rV��,y� �vc�F��y�g�AU�ʨ+˵@�	il�CW<���9;��/�*�z 2��SH��p �u�7nxp[	�| �\q���d���z�a ���I;��� ����-۽ l8ߔ�3X
W�94� <�=�S�Ctk�Z<�%��΀�1|� �?�w�?ǀ�
g�Q�� �p��"`�� �?�C�=��Q} w��]3 �-_�|b� ߆�}s�	 Q*4������m �YyF� ���C{)��ע@����� X��g� ��P3]���nM��`�L���`2%�� 5,�~<�\�_:� L_Z��zh�@��!�= ����e�T��\L�� (o�ݰ�~R�$&�	��h��rw�Q~f 7��K�H+D�� ������7�a[p��q�S� �h��� M{ߣk��;�Џ&�����Nos�T"��ڀ�p���,� �+�� ������A�q>�c���@�\w,$t\ >ʍ�j9��X��,
�`0�Q���������W�.tB>�:��8bȏ����7;��x�@��=z\2�S�U@_#����˟r�:��~�`VfJ�{  Sw8-����X�@��12�� D�T�H:	ۀ��T|t_ s���`�/`���K �	D�l� �zJ�#t����{��0- �9j�����Al���`s� ������C ��Q���:�;1H��`0� |es�'>{S ���@��Ә.ҋHD�y���0¶ ��w��L����5{W\0@�J�s� 6=͓M?a�� S�!�bT�� �)�cC� �4�35 ^1=����4|�� G��8$ �;_�X��I��q��/��� �],��gYrK��-%;"�
�'JZ� ��N��`�[�w���C1 �=b�G�+ 0/a�W�6L��x8Y 0��ʟmO �[@EF��=�|=q�p�B<��V�8/E��z��� ��)R-�fX9��2x�`��� �v̴���� [Ï8~��Z�n�K�܉%/ ��d�pϠ8�� &xFgٹ��� I�Z@X�N� ��l�˽� �"�u��� 
�e~U��� �Oh��1� ���+��xS A�-k]ؒy�!��𬀎r�� �9)hD_��y�L!qK�)M���� 3\u"v���� (/�X�` �]��Y�a�{�UO!�[M�PyŸ ΢7NL5
��;�2 ��ʠ� �����65Ԯ���) ��L:y�K `�Y��U2�	��p��Hx� rI5z�ی� ���;�Y= ?�l)� ݚ��+�F� v=�@ъ�W~��@U���Q�@��s^�	����3ͤ ��[���ur�Px��I R� ��#E3�R; y�m��L�M ��A�>�� 2�k�v�N |�4�!8` �,�w���Mb���AC�Jp G��"�	 �# qu��=����`�����"���t��<�} ~��� ����Z�"� �� l��~�CKz��`-�; ���$v�� �D��� ��.7���;Gs� 6�a�ۤ��^�K'�A)$�rʽfZ��.��u��̓ �$�%V�G_���>Y����'�~LfO�!�',��l�k"�@.m��L�ݙ�?���Y�����vKå����<�ܿ� nɳ3.x� �Q��f$�7�� �x�Evz ���������`}�[�w �WV~�KIg!FUp��v(F� ��XEYu�+ �{�H��|���8s ���l�i�7����p�NQP� � �ĝ�~�"�t 6�-0��$f�y ��/Y��o0�Ъ�(SM� (�~�`�z�  _���#W�v� =O�Z߾X�� ��^��.�?���*�{����GT�m��/7�� p���� 	L-�O�] e"R�S ~+����,� �(�����G5˰H��] �4�Һ���"b��9�Ł�S8� �� J�,Ѫ n��+}�|.i ���%(�L�)Tc1�7���{� �,�(AI��,N4  ��
��x= n�	����< u���阐$ ?��&�x6���;�d�&��� q�ބmB~ 2����K]{F�S.�0�F��0�8�������k���,�u�c זB�#� Pį�n� u^-�;)*� �wB�D��' �Nd���:�ՠA������o� �7(� ���p�j;�� �>:^؃ '*���,�! �;�ʷ�x�0������Z �s
�;g �q+�?�֌^�'/G }~|+�� %�L ��\�5V 4Z6ᗴ� T�r(9���C/�s4�y� �Z�dx�� �j/�N�L �@V�n�v� RT"�c8� ��`�)2j�Uڮ�pp�3Ic�Ԭ���L�m�] �|U�	� �I�o>td� ��D�@�k v
08��V�,uw _�hameG�>�3����x� 2wc���� (���]� �����V��</ڇY4oCa,���G |�~���� ���@w��b�^v``�Mi�߬�@o�]B� ĚȾ	�~FƘn�1��H)Á�S#��߅���u�W�~, �'�E���B�p�g �4V�w� �D���,(`�Þ
` R*�e��ʭ��]��,4r�{���V ��G�u��=À�28UBR�\�� X^�w� WI9�o1�� �x����k:V��nb���o�N��`���t}��E0c�� ,��Ø�0mQ������-4sոL7���z v�U��cvx �r*��As_��q�X� �id�\5��z�":�0���ȧy ?$�g9��R&�\Z �t�.m 5ԩH&�`4���A��p��� ,�%P򧶗�V<Y2 ���� Wr���:���� ]�V�Q ���M��% ~;/xVI���C ���7B m;D]!�� Q���@�>F ��_Kl;�] �{��Ϸ�|5Xv= �>�l������ 4��D������Sf0�K �Eqж�$� `�(&R_�:<����e�7G�O�@3k2�,�>)˿����O �{���C���l�3�2 =�O����� �8ذ�J��(Ż� D%.q�O `�861\2A '��X��F�cT��_�6 �»hUG�4 �)u53��&^� އˉ� nP�m�/����I�N�#�j9�%��oL�?<�ۊ� f9�A��� u���wНv/~<`*��m�'��k����Q�E�둈g F&��\@S�Me,��~Z�8�;	���1�.��護���kl%(BG ���z t�y� ���&5�m �u�h�sܫ&� �� 8�����o�P:�� W�I᣼ ��$��X}007�WH:������@�Ș� ��)S�{�� �8u&�Q��>t ���x}J~; C诈jZ���VǡE����K�9��I.���n��&݄�5��w���ҕ 
27��*gv �ܜ���1�r�@r> ���穭<��vZz� F��}]��Y|�j�G�V���� ;�M�9H�*�ׯ��S�Bjy��.������ ~��ȡwn X(��k5u �\�~��3 ����(s��=0�����C+ �\����� ֖e���|?� �-�������P�HQ' ^2��Vz:�Y��Jd��& D�H`���S�,�T��0}N��/ȨA��7���)�{���1����G�&9�lZ����'�a�%��tN�mL;�� �R�	�] �Z$Ca~=��e*�1��� X
���5�~� �,��"� �}�5h�G
p�;���E�� � U�)�n��� _���S��� ;�+"<��~ ퟣaX��� prm��ѕ�˰��sI9^� a U[�E dK��Q�� n^�����7MZ�Ӏ����tC?,'S@���tF|*s���XG z��� ��Pm��� *\w��O�k� �+<[&�� r��.��*ѐL �#?�G7URH�� ��J���@%S	,5 Y�O��:� ���v6d� ��:;	��0�
~�S��UFg�����|��2�ѮCа0%��ߕ���rvF0�A"+ȗ@(��><����c`�ʼ�;wΐ	/ �Uˌ�B��K �)��7iE 0�����o �1�"�s�����JW�� tؔ�ٷ�� �@��ޝ��[�B�
.� �p��;{ 5 ��#���9�y� �z�`��Y;�� a��g��t 4k�J&ƿ ����{:�J��� KL������ �p�m~�p�� ���2�� ����w�o� ��'m,V�8+>�;h n뤈��f X	ui�+�j�4���� ="�����H�۳� :r�F �C����f6���>��F��E��p\�,w! �-�D�θ�X�� M�Bc[0/�� ]b���V�����{A k$�= �/�q'\ �OP��
f䄳��S !���˸#�xU�䠘E�Gp n�]��#Z�9N� �We��x ��f�H�	 o��Ci��� �AwmU'��\�{ %�-�j�B�J�g�I`�zy� M���G^���uށ����t��#�xwA��r� :h-f}�� >+o��B��e��X{��f� =����\��I� D�ɏ����i�K�+ �_o�驚">����Cd xzZ%�:��h����1L@��p���Q�߁�����& �F��m#�o �v� 6c�ٔ�=m�gU���� ��ɾ�)?=���T��/�R�v +��ڬ�� V�*������
���kn�٤m� O�]����x�6�j��> o����������t@��ȞD L
���;X|���J:�v K^�l�u,����D�pQ�,5U� �C�+ּ ��͒���5�B��D�z�ؚ+� � I�%��*�Kj�LcSOHW k/0��'����9Ճ J�N�H��冕�F�4�V� }9�t� Rm��"j�]
p8��J���{���	 Ǖ�&�\,� Ɨ�ϟ�( ��f���D !�~8��p�����^?A�
�Jw$�V� ��kʧW� ��%ޣ�Q ��TA:y�8�s<�K����G}=7��$��͚ŝ� Jn,�{�6 ڏR��>i [�J�c]��;���˧�@�9��(�����u ���� g�>GN*�{ �s��3Cc�
 ��R���% h���_O�* A�J�Q8!�����V�>�j�^� q.,������5!�`^�r� ������ �F|��d1 wf�ʖ�^@Bl�8yQЙ� �r�
� �6$GC�t� hd�Z��U����!�[��jN��`�|� e;�M���*&��v����p��� ׯH�6�`F ��J������Q�A���� D��.����o�b������ ����j�X-�+�n��d��Z� �r�M�?�"�ס�#4�a�~��� ��|NlD& �ڶi}ݰz4 �?��t �D���#8ҕ��'��������`w���W��r�{>.�ީ�ˁ��Ip;l `#�z	\)��� ��?h(� �j��%���O܀+���m"�O���`��I��# �{ �Y��Xn߷u� yNFkְ T���), ���	f�%y��Nҍae�� �����?0 �eΤ��1h������� ��ͥT1Q�G	[=�xdڊ��P� e�0�Z� ��2���� A������ ��2�Z�e�� ���Rg�p�,Q�� 6�����@�=�T� �@�����-η鰣q�
v8 :�v����$xXb��=ah�Y�/oP� ��MS��0;�1�� �h�-?|��Y J�<W��GCQ-� ��7)5��|���`���F, bY�ɣP:�� ���ؿZ�? +�Ģ�(�d�r�:ۀ4�� ��OM�~����&� �RIZ T�C����s�>J��7�#�W�HK�t����x�T���!��,/Ǔ�`JAcg" E�ꔑN�< ���,�3�yo��|�L ���V;3�7k��p���.*(��!
��@�%�g�s ��w�6^ ��ĉn%�p� ����1� v�CADt`Vyn�"���F�� ۝8ַ=�� ������� ��-l1@8��p�c 7�zW�0F�JyI |�>�q��#W���� �95� >��b�V �|TF�hX�<� �s�"ܝ$ #���.`�:�����:�9��i0��<��8`��Fb�g~uH�l}X�P��4 �.0����v��<1�E��:e Y�F���� m|;J����8SNߪ �����_0K�>�=��A���:o2���ܵncN=q��b����e v~���8�� ��mr'#�}� @69�l���$C=� =��1�� -�"��Lפ�p��O��#? ���(�;ݦ =7��gdHL`�`��0��x4=� �zGW�*In ^o���#(m>T �F$y�?���8�}LpR� lF)%�@�X�e���*���� �ix�z2�%�fH&�Y� �	�/|+ �J����[L��@�) 9�XB� ( L��T�-� ���@�V� r8&�I�� ̋C��Xa ^��\��Ӹj��)clË��Fy ����*	zm�&��l c�� ;��`�!Z�m8*�vb�G��eǌ+TM���IHA��^������B+> P=�ɫ�eF ��,� 2��S�� '��/�Kg�a ������(� y�I�k ^ �H�K�2>� �v�'-�r��zO}� mA���k� q�eT� �p����(��������&$��$hi�ޚ P��^�"��H5�@��A��	8ダܸ���:� ��}5�-{01d�i���6(��#i4��9� ��T8H�2� ��qV3A�*�܀ ��'���U�|p�m6L���(Fģ>V���}��� zD���E7� -U�t��<a z��@ �esC(�� "��A�x� �\L�7m@b r�;�:�T"��������<9�}x� �4��)d �����ũ�Ȅb�H��$��:D�/�g�J�NM i�l����@����At``��`5e��� '����m�	n��� �`��W���f������ ���+�9 ��q'Q�T~ kR�y�^n�������|Hlj� �a�v�U /����KF��G�?��t� 2.��yl��@��Pt�:��gU� �۵�a�6`�(�wY�b��= �d��.�|��\p� u4�}�2+,5 ��iK �� ƹ3���P�������� #f]k�/"�6��x� Z�.����`��nX�A �}�6�	PM� G�ԅ��J�kF�и;P�}xu� #�Uq�9k�e�\��O��x>o`{�J�� �3(�%���:e��A�j�
� ͏7�ׁ�	��<9`r7��E�������L9p	tc���-p�� ��"���f�8$�OW*H�aqS�I�߁�4�Kt�| o*�:�9XXۅD��/��Q@��_ 8IG#�o�2��|�C�F���� r���� ��aƫ�* �y�����Pf�� �k9[�Hհ ����J� &#��%�	B|����N�^�b mI�}j��'f�vd@�~a. ����!1}[��σ8V���Գ�X1Ӊ��plϱ�������_D�{�a��R�A~��� ���� h; ��p����b�NG�@=�����U� Ȓ�2O�`�-tŇ#:� 5����� �
��1��> �O߿�ٴa ��iЄ}Y\��hs�рf�] �I���0�;ª�r�^��,�� v�,9�'�� �K��&� �g��nq9�ƀ����|u0��U��y�Ÿ`�ȀퟟЂ �N�� ��\�oA	�sP� T<ܢ
�a�����&��|vh@O�"x;�	E�8$�I�ذ��Yt��wv@V`��I� c��N�6 ���+)��  Iy�*/�qlNk�h��Q
�s�T�^$jy 0��R�(��I5	����� ���~��O ���U� �6�F�L�<ɀ]p�[�*QP�� _���� �>�*A^	1�um�s��Ū��8�ۃ� ��B�$6�{�� ���+1߷4�IAeLV^j�� $Z�v>�AM g��/��'}�?|�5�� 4���g�
@L�+��� �WZ��&�����j�y�Ϝ㮖��>�2p�[M'u<!���7p���k�����O�|� ���x�  �*�? ���&m_ (H%ΪL�[�������������:jk� ���ۊ�8's��� ǈ���/	@��9d� ؠ�IX�� �� q�W� ���zh-Ev<�#�>��d+�.s]�L��=T�����v��tp��g��J� -�/�L��q�v_$>�π��E� 2P~�;}�  ����<z���#� �K��b�� �8���T3�J����40 ��D=r��s��[ yRK���P �¦*��g�!T��P�>�� �|lܖ��>h� �K�ב.��a�)��#F�$�� l&+�1���#i��`�1=��t!���p���v�Z�����x����c���Z�P�
����� ��� Ӄ�.��� �袉��2 K����;�P�0�2-!� ���;f ~Մ!��
�B� E�R���\��x������;�� ݹGP3� �q�>O��� 9�	�N�?�d���W��}g G�%a��3J oP�R�  l��a`�x�1� �7���+� �Λ��%����-�.�L� ���,�� ^`T����<>�� ��y�b��~Oz������Q�� �S|X�Jh��|�d3�Z������ ����P��* �U6����	$�π�r�?T�xc���\y�9L �O?Ǫ� ����+��' o,��-��6����� 5���1 ��
L� 2�U���8z�+ ���`�r� j_&�w� ]����`�����`��b&X m=qYN��'hg0�����hd� 6�?qܻ��ND@\�E���X�Ɂ����C ��W�1�;AP/l�M�@�F�yD�n�M[�\9P(fX��Jq:�
�A�����H�{��HёR�� >�I@�ToZ&{�Հ�w?/ߡu'�~�@�HYCoj,� ����;w�x� �^����p�M4�߁#>D��k�=t`�x��E)�H����������YQ�2Nx �����7�D ���eX y<@u��$	G�� Tn-V zi,J�=�:l���|�� �,��J�p y`��MH������.y\�`����f�"q�jU0�2>w����Zf>q���zX1� �rN�t�	������-"�@<f�t; ���������$�Հ}�-��.�B�		ԃ D��7�p� ����fgE -�9���^�;�8:�Ļ �J9�R{��M�����������vn
�u�Y�Uz �Q��܍RN�ҡ�AB0���M��^ ���1t2 �`���?���}R�o�6�+� &@������F����_]�� �G
*�Ih� 1mS��: �������>0�-)o"� �t��4���H?@_e[��,�0������M&�.��_2 �RoS)h����]$����� [�9��W�&Ӫ�:�-���px�F#�N�jx9 ���l� ަ�/U
g� >b���ld %�@�7� ����K�͵�QI��N�C��/� XAoD� ;=��Buy3pFY�!�( ����u�X�3M�`�1�ڨ� {�(��ҭ� l+C},�F t�wW3SHTFcorH��G ���3��#I����� ��Q���B�`�AO��
�d ������� \���; ��s�8[r�}�`A�t�&D�0&��5 B�+����럠���$� [�K��|L}���cl��{0ЀaU� o�3�� ~� ��s�?�0����-����"�}���! �?�`�~��������t����| �패ͅqG �����	� %� ��� �2M������k���h� 	�`�(����1ێb�Ԑ&� \4Md�|� ���<m��� 0��&� ]x軓ZU �C��	�����C���꛹���)��D\9��}�'����g��j����� �E
A�uԧ�9W��~Lv1 n.�ğC*9�Ѱ 	,�o�X�q�Br� �G��]5VLDv���UR���哷��1���� Bv��=8��W�i^"zQ�����!霕��9������ g���Q�z֧n��s��xJÑ�>0�v��\<� 1%���H|F�8	�lRQLm�Ā���$HezI� ���� ������P�K@�!
���3�\�� �a$�=H��>��!ZuTH7 ���4i�K�&�}���l�y ��`ݛYI8 B�Q�> "��L��H�M �Z2��� �#�"�T�QJ�+� ȸ�� �B����0pX��O?;_`���- "@����� W�F��+� �EA%��� R	�C��|vG ��b[� �0iߪ���n�^B5n�<��VE4� �W��a|3=�x~c���iE e.w���� ��	��'\ >-p<aԬ��i���@�F3�8P����k� �VYR%x� ���'pδ�D�,e�Z0h�.�+�˽0� ~� vr�2���� ��I�ē��Q0g�{�nk���l�@��HP��A ՋLD*:�m ��ٍJ�0� uj
Y��������h ��b���c� ņf޽
/ �sY,��#���|o����^�=aB��w,� NG(�z/mf!��p'c@3��0ZA���{��h6�d��0�����'�M�-��HDG��g���j��L8 ~�G>��%���w|�����zHg��a �2 �un@��q6(
%,P*L4� m��c8�'޲�x ��6 �:�S4� �%���~� ���5Gcfz��oa� �B�u���h#��l�oH@��5�7!bd������ep�J4�0 ��am^v� ��dbL]��% �9�����X�#q��K[�ebg�j�	3!+s�2_�&�M8�к$ ����Y{���y�� ���/!��k"�A�}������#�Ϊ�g̕�����~`n�q#H<1`f�?����4\-(~� /'�^�v	������`6n���&g�!t	�7N�H�}��(`q1?�@�7*�| 4X�#�������S�s/=Nk��� i��4�A 7nHKJC�}���	$��HYv
m�>����fR ��vG�4, �
Bza�� n��W��� �>�I�@� %+�Zy�˶�2��^3��1�W� ;��4V+� �1Q�-�h�?v�p�u ʤ��E�p� ��7���˪� dϔxyO �^��,j� ����3`�᝛d� C0P�{?Qo ��"�l�9�L�vC1�Z�	���� ��>��S��|� ��Q2�a� �Nژ~3�`�M9�b= (��Z�4p�t��:�X��� ����zO� 4�f����51�� ��3��e ����9J�v*u@��`2��,����dyq� h�7Y��R �򷻳�� ,�å�8h ~�D��u4=�@-�x� t0�<?�* ����(�A��s'�E� �U$��)%� Ǝc��!�`+�.�z� s�_�b�W��EȲ=�yE����%��S�A��'��O�*����@ю`@"|?���1P5MUt F/j� +�
�,^� k=�%��=� (��[h��<,��T�*��݌�:��C��i �~����Z 4��sU<@	�S�'|��R�pM #2YO]�X �Ŕ$� Q�?�}&0� G3�X���KE`�W
��&��\0�'$� �:/W���bxa&�I�N�tY����������@��� �W>6Q�r���/�t�.� ��7�f�Q� !RC�ܙ� }9�˻��%7ٔ jᴍ�� saZ���`lRݏ�����s� {���^Gv� �F�zA��=��iߒ
$� }޺O� ��z�~o �ٝLg�]9�� ��f�yL+��g$�u�H{D�<���j*������ �9�`� �~��M���%�}�񒀈�R9�T�|@gm�>� 1�jD7��y zi�J:=d�F��@�\]�,�~
�x�g�p�ڔ� ��*F��o�c� �S/klKX ��3Fq�(Z ���H~�GR1W A����H0>n�2)9�Y ����i  ?�ȸ�՞c���@0�b��s�-��Q ۭ$)�ƕm�:���	@�s(b��6�V[\ �X#Z:N�� O�G���w_$x�� ���{8��)����* �a7j	L�b���
�ڪM;��/���5p��|� t�V`kۮ���@A=��p ��~}��s 6!�c$z �⽧~Ýa�r �X���(���=�_��go����� ��|Dq��� I��UZ$� 7xP�_W�� Co	4"ؾ|9��N�0i )�H
1� ��{a��SAįBm����$� 9����%� sz���!�I 8�iyC�����σgK�ت?� �c�zP��Ǿ�����Tl ͽ��ڗV| I��LM��*�#�m9� �眆��B�q28�X��\��WC�$��lDj�hPʅ��b�ؼz��#f�
<�eA��������?] � ;i8�!+5 T��f�]A 2h�a�>�xBM*q;dA��q�� K1��n=sf\�WC��� 5��Ɗ� p2  !`L3�� ��*�yA�u�N�L�����`�?�1jK$Pw�[�. �,����\��Y3�WiL�����q;]��1��'��?�s�-8tt=:D;��` .�u�t<�� �*�
+��32҄�����������/aӱ��C/��w-��5�#| �^i�o�D`qb �c��/ #�\�6�o �0�羋 򮫄b�h� ~�)�+ Rc �F���p� ����U�q �A�-va�X�HW�V�'�h0�"�=��$5�o �U '|�.�H-@�d����p�y�?/�G% ����Q�� w�~�{�� 4�.�d�iE�q� ���/� X9r���ا RE]3��޵�[P�) z�о�ɰpI�7]��3d)��8���žp��;˙ �0�G�* �`O��v�s	���t{��n �@��G��|>�� �p��h� ,401��"9��=��*6�� �B�7��_ HY�S�~�� ��IVPٍ�>�+�L�o�x$���a�@�'�(� �)��n�� ?��Jx^��H4Z�D���n��w�A@�bc���S� 8!�#  ���5�� c�R'Z{� D��%Uz�?��"[0 E�X�0�81Ww���hxR<�:wa=;��9~���o�� C/F"���<��6�T�qL 
���c�2";d%�0R��:�0�Y2��>�!�/{��I�.��Ǫ�GD1w΁�&�#��;��_<q�@��*8�����!� ��P��F ��X��5��-*@�
6؃� %o{�n�� ׼�?:c� ����+9�0�Ґ&_8,�?Q �]��= ���%[����|g�Ҟ��9{h�՟I� m�]�rC ��f�G��u"����`p ��%�ܪ�� ���1���'�Aq���*z2�7 ��n�< �5�{Hg�? %��s�}4� ���"\S� -�![THC k�=�f�1Ypz_ ��$AH� -yص����f �l:�W's�8,d�ŋ_�-j�� ~G���2�LR�f�
� 	ADWma`6r� Ȩ�0��"o;O9ր<&YW6)�`7��r���8�X	T��~G�ȍ
��HO� �q?Y�1��� �Fl��]E �b�e��� 0�Ǐ�t 
�+ J����2@㨓��0_ <f\F|Ex~ �#�z��� �*�Я [듔ј��"������7 K�L>S0m�xe_�(��`k�`�H�/*��a����$��6�M�|,��&��s+�ad�.��f{ g��>1������v�����@�L���X/cװ�TbaBW�Op&�lN�p�w��3+�=ـ��)��=3ǉ1�J_ ���2��!�%V�L �.�B��e��QT��@m��	 �U|&֬ ��ƪ��� ���c`="���N� ��L�a�*���h���P��@� :18�OR>���t�Ur��i�0g�=�j�~|`�-�'r?��K���V����#AL[�2���X ����g�^��� ��5��jk(�D��tz>/0��i��@g�I~� �_��Y{� ���gn�RLp ����ǐ����<�߁�7�(de ���������z�i�:R�0x� 7��$qZ8>�%T��f�*�Y����C��������d�� ��b�r�;�X:/H`�}T M�Wݓ�<�Ja�+�� �-� �����{ ����iwx� X��92��t1�!�'��[� �����c�?�y ~�g�I�_� ��B�.�&[o���P8��� ���{S] ڰ4Ϧ9 �$3%p ��w~�8�ne��"�v������/�f��# ��[�� �?�gH��@��JE�Ѝ,>~l���O) 1�WS=� x+���X� �*y`fo Mm����� ��8p�A#��:/Rr�ܪN��C�����|?`�X���.�O� ]v�HU�.dN�b��KD�� Q)V�A��- �S��``�A�F7'ZV;9� �� �W�x��� �i_+�5�?͆�h����@<�_�=CJ��|�z� �>��G�� K%�tJ��[:�-'D�>����� N��i8�x� 3�=���5� ��o����������u+`9! HlG&�M T���ܓ#1� `F�"eD��!&P�;��_���P� �ȝ��� i���3�km���0��5r ?s��`7��H��2��Zճ ��y9ͨ� e� ���1;t��qX�� s�i�Bu�}�W���������=G�,g��ϯ�vn �c�� 5�A�4�1�@�̓�L��@�A �s�w�b�@ iՓ��k�U�3�V�;�w'<�^@ �9YA�o� 1�	C �?��=�]ޙ�u��� G�_�A�s%�`�r& ���Q���J���p��<� ��T�s� �2���B�� <�{�W� ��Z�6$���;�3��X&: �^Ӡ�ע����m9�� X��O��]3 ̆"�P'R� z$�h^(?�P<�g bG���@�c��?�(����� �y/d��B �]	b�� S�:JX�*��wj|�dۃF���4/ @'��8 ��X_��  �"��o`!� O	Dh�@Ɇ����d4����I���m��0}G�e�pШ87k��J���� ���/�w-�07 p1ʩ���K}�g����B �	 �������@Fq �. �>�jR	�=��|4�����tgJW��0!pC(���m#�r��/ 
�ׯ��M8�� ­e�f!�� )�K�+�hsl:����Y�����}������J�hX R4���( 0 ��%Oݹ ������P# �����k�� �V�w/Z�' џ��5Ri�� 6�3�W��yt 5����p$�u��y �5M(� gQB�Ok� fP_�Hh��� �IW@�1SM�0��`t�x�3�b��S���M�� ����t��|�[w�9I��}��\��]�H�e ���d�<��@�.Q��� ��l�[?���^��ΆC� ���	w�XfnC�'��a �@�ߛ�̦w�nh��d��\ B��[�A� �;,�M�λ �p	)�:����@�th���T����@�~0�u �4#�;����`\"�ߌ 	`�!�h"�$>��H� �G; ������9:�2\��� ��Q�l�Yf�#! ��2��;�a�� �w������E���Ҳp;�ߠ��X��p �Ⱥ���ɟ@��$ N�Jⱛ�}� ���&��	�T �(��V Ͽ�^<�n� Kӧ[3�so QҠ@G�R��
@�:�V�i�N1=l����qB�?� ��(����9�<����p�� �،�$e� ZJ�|%� D��޻0�@�����|�{.��8��?���<�-$�5�$M|S�/�ۺ ��ao��� ���L�pa 8>�
b��tD���"��a��q|��6Q.5@UT��o���\�P �2슨~ �U�T$���*"@8jZ�Q�ȅ�8s{��\����y P捄bHt5��`���J������!��E�_��o��i%�U�p`V���=�� �GbR!8��$� ���4H� ��Ù8.�P����͟ �Y�H>�z��;M*�
D��V�W��p�K">�-�����_��N�x@��@� ��ɥ}�!h�75�Ӱj ?��zB|y�+>�0�G;Ž�Uǧ'\��8�P�� `�D��-�¢�M�1 ^�BC����	� �i�o�E!^�G'9�|���l�J|$ �&ᤍ<���f ep��U�Йa ��tzZy6f�$� ^*�) ��|Z}�b �q�̒���r�x����B;�8t��>*
n��=��8c� 4(��� �A�5hK�@=pf�Q��d�J��LC@���:�s�a�
IxT� ��Z�rQF ��э�|�� ��^���Ͻ hӥu���Þ
�Ԗ:�m�[����J�����|�(Z� ��rsM�w(7!����,"� L�X�� ������r��WʂL� ��`������wЀr���i�n~� ��߇ cvb:��fa>A� �C�pW=��O޴����{���k�h|��X$(�Ѩ>T��	М�@� � �oC�\{ m�e�qA*x�� ����J`���!�6 ��"�x 	��4ڇ>z1 �?S�ކ�[�F���ܐ���ʼ ~�
��zS}w��%�f�|�T �a�U��� �0��!�p �,�}��`y(��bs� ���0��j��g�[ #�M��o�VF��Z\Y�T ��r����y`8����=�}����e�>� �K9.֖E |Y�W���������ͫʙ@ ��Ǩ/%t� �|��2�֚9��s��0���Kl����p��y� ��@�2���
�:�V�S? T �]�	��F�e�j���,��z �M��%�� ��(:�]�|!+w3�v��I��	�^	�d�P�R�O� 	�k� ��wBh�� *��r�>�% ৈ�h����yk�5��, ��C���] ��=����� ���K�2� 8�IS��� OY��x4�:T�$L l�Bo0���e��|@�: ���7���M��m`2��� �lP��S��Q4P�AF��C඘���r�c,���)؁?9T���� ����D�VG��� �k	�ig ����I(�/ ��,�	�y� �r7qW��i�Y-<��,����ȝ?N� :/��� �D���?�$��n9�Q��� ]�����$�&@ 1�Qn�h :� ���� qpN��Z)�8n�QP��F�>	$�MK�����8 =��t���,<Y�l0E9�� �I*�L.��gfv�	Ġ����@a��}%�:����
n=�e���1h	 �_���bv�Vd/���� Qp�T��5@ �0D��,� 8�����>	.
�O ��K��z�X��9I ���2�ʹ �ZoB�~���,�L@����I!��_� ��U�:
F�"��]��*�fS���x���!=��t��p�����X~�p]cC0ˠ������"��ТT+���U E����8��_9(�!��f� �yjut��=sv��>ۦ�0���������`��}�u� �4YA<w��+��$����'�O?�*��{ P.�/Cx�' ����d�� �ؿ��tE�W�Ȱl�� ��#��'UxP f�B9塗_ |����Ө� ���59�7 j��և �B^<f�PX�@9;��� ��,>q�g@!(��n��"吿 ����� e� l�(5bxm W�|,�]P�!�&��� �Z�-�� ��P�"�8�V��ć������@�� �إ���B���84�� a����,`�����up�* Ύ��y�s�Ǆ�W�༥Ă �m�q��A��j=.�A,���2���^>�Z�$}��* j7��̈{����0�I�lu�����c�� �X�TH�:�<�`mKA+�5p#C ��{���N�dx������� 4��圇 ؞pW����x{�	n��$��h�{� ��F$��@a.C�&�v�"�8ME �Gcg�5&�u�T��%+=ǸЈ� {�@7t�" U/�ge%��q4CwD��-����	�{ż���W )��U�v��_�=we���zX ����ck(����Y�-܁2 �� $�:�7	�����(����.��1!մxX���xnt+ �p�J`���f6U�0ʾ�Ր��V����a�m��)6� ������ �_����X��� kV� �8��zf��)!��W/ ��F<%	 ��&�5�s�R���{[�ZAHֺ �5�t�_:��lL�O@|� � �ڸ��}���d�|M` )� �S[Z�~�l��#�e����	
�D ����?#���x�(9 �^��l+d0����%����@D5Y�4Y*����]�WU�n�6���X���r���"��䔌���N �T�8�q]�.m�r�z��h <��K�uL =��I?��Q��s ��~��"��b+��"�	�wH)����K��h�%��]mi� �*�±܌� �ُ�jݎN U�뉜-�Ӱ���\�|l��il2���v�:W� g��?��f�� ?��c�����*�O-୫�����"�p�. %�b�_�w���-�o��xF3 ����l p�t�j��`�(��A9���xKG�J�� H�}B"��DMy������%��"����� �Zs�q��{7}�P��������c�������)�pۮ�� F��2釞6 �z�5�Z?�\�C>$�������@a���{` C���k�f� ,aA=L���@��يsr$`o��2��<!閄�h�(,��ϺX�	�} ��v� �$V7ujYH�M�l� �y�W��Tν�eQ�q`p|D �a����ҹ���gM�����e� rv�30���9�M��LF����iYag�@q��=~�bb>h��,�*�?-(�4���Ly�����*��X�x GV�a��bZ:ܷ2����f�*�PT<D��]@{Ω$ 
�EК�� �蘐��^� �\h��UH,�`��Ey�`'���{���ٺd�x���ƍ��?�]�A�S��hd�>;΅?��^ɇ� 0b���M'�@ �y�D10#��x琌n'��`2K�O ���M���x h�.�"��*��m%�9�^BK���� �" <�g$��, ��p���J Z����l� I����Fy �Ӕ �2zc��⺵�М�yM�~8�	+����Q�Z��i���)�����W�,�=�Fn5�>R[}��B���E�����" ��yHD�@:I�z����3� L�w8%�R[QX � &����vU���a Is���ʆ� ��c�wk� M�S�Hi
������\"f�@L��Kw�� {�'� CAڹ��q<�m�%O����e� ���雦M]q��PpT�)DQ�g�|�q���,���$�.� B�|1IΌa��I��:��o�{$T '��v��ot'�\$���ܦ�	{tw��,G�@�vN �ż�5����Á �o�����@pDt��]S��p6<,Yz� �]+����Dt\h'��&7h ��[��C}��p@�a�˱0�U O+�zQT4 ��ͳ�� {��B=3�, ��LI�4�^}� �|�o�]��$"A��� *D�~$Y�uQH�|�ht*��B8�����������
���؈�X l��s*��'(�1̏��� �-M���T �XWYsx	� 2P���� 3/�]7�t^����+@TL�,e���������D��Z>��H��h����T��<���8/ �C+�\3�i�ߛZ@��Voz]�NY��1��v���T
5 ��S�Hd-�t�*��&�Ӹ&��<�� /�3�$	�s <��:��?ؼ AʣKk�E O�@��,f�X��� ��IH�����= �� T�� �����1>t �a`At�< 1e��}�F15Ű�Y_9� ��$5�my~6Q}p49����"��u�k�+ fX��y'���?< {$���G`8h�l����kH�  ��Ȫqo=���S�^{P*�q9��ﾂ~��m���C�y LĶ�;/���)�W�@�J>�t; (���%��t' C�	��w 4?�R��~ �"�c}3�qh��� ��G���QC�̌�H_˨�,�� ��+��5@�yZ�����PU7��%�`����|�r� UB�`�+�y� >�!��pr D"�P�GV �e�_��Pf���:� 0`�|�� R��Z�U	Þ����0V�6(�'�E>?�\�+B�jcz �-�n
�s�N@E��ѭ��g�)�<l;���>⸀M�D1B�;��t�R� l�XNɇ1�,�zqդ�aH� &�ݲ��<�%�r�T�ی Ѱ�'�Z� �8���h��3����s����:����-bVļU�5���TF�D{iM�� ���ڷ�в�. �_���Cqk�mr��8���fB��X����/k�&s; ~�z�vxT��{M�������`�O -ǣy7����JX�$���0�NKcT�|�
&����� NҠ=��| `p���{�/���� �G%̨�[�ٻ�Mଈ`�_��h⠔�yK�~ ��p����:�� �	IGME =�}m����X� �&Էl�~�5ڄ�v~6 �ɬ?��f	�zi�acs 8�E��XT7@Ѣ�|$� tdH`oۦ	\ @ ޵7���3Ԩ�w�,� ?�{&�oh� ��b7��m ���ꁆ�:��P���%�@P���#���4��p�	fP0���}��
gu��>�i����q�è���́9P�u����
9�� o!�������K'�)�̀\ݪh�A�P/�'ҳ�X���l����X� ɩ,خ�;��R�F����{nJag�/�A
����F��0�0��E��J���`d��� �W>%�O�S3	���9�� ���2}���$M� ��9~8�+ �W��p� �`�s�A��ecf�7_�j&p�t|���7�� ��(���9�L( }A2�Oکc���='xw�?�� j5>8dw`A$_?� 4ֆ.\O%�� �T��u�9� �I�N[: 	�2PRU��'��Mf����c�0�:�L �o���Z�� U.�I%� ;r~F/!�|�wy)�d���s� |'Z8?�r$�9���B��k�j�	�0H�bS�q�N�̟� x�u�>ڂ�����l���v�Voc�ܭ( �J�D�i����Y��L R�T2 �"S�O� �p�/��:�e����ÀaV�~d�m��'��!�0iV� C�7�R@;W �F�p�S� ^�~̭�Ŋ#�) �¾�28��$G� �O��L\) J��i2��� ��c�p\��;ߨ�Y ��DQ�Ls=.zQ �, �Y�CQ����b]&Ỉ �p~���{�7�� 8ف�� ��h�w޴�x����T��bX��}���_��,OB��	d#zX�8��a&_N� m�H�����.���@lݍ�q�;���|g@ɸ96� �45��`���܂��Ր�|��m$�E<`���A?�0 �1�O$
� �В�)	�Nc�X��!�2��1�Ԕ m�d�� 9#���,� �L�)'���J��� }`\�ރ�N؋I<���� �&<����o�@�h��1U����zXe�{* �t����	B�+�t�"�u�t��Z�f��O�Nx�
&�h� ��K}��� �b����n �P�k(S�{b\�8P�:>�ҝiy�Cq�v������]�5X<�u�����
K��ǼA��Ц[ 
`;s���t'$�� �k��l� #Xv<am���z��)�����!d��_�0x��ϯ��b :���&
e=an0@��$F�"�Y��&7x��;�잨�
\� �ѽ��<��㑾��T��F��S��?�q+� �y<�f�0�Z�̂aS B�Ҡ�@vfrq��'p�Q@���;�Py���%ۇk�]>:[�0�!A� ��@+�qv$�~���b��Az�Mث��3�CL !�r�`���*���F��g�2@�@�?v G�T�F�k�<2�w$��< Gno��Q�0ԑjRX$q���%�D�``� ��� ��wv�i
���
T�J�'ۉ[C�"� �s4����6C����k���Zh�)ۋķ@}1۠�j*+�Hz��@'q����p`l��}�@��C"t)O�p�f���!^K"�
 !k��>��A�*n�Ġ�g��]$��s���,�΄tK`&ۊ##� |ۿ�< �vt�����^���L��f��F�M"zt? XU"�	]��;\\&����
��`t�H� p+����u�� ����f2��8(Q�o��r茵����%L�� $w���y��x��xaS�� ��)PK%�M���FB��z���(��"�I0$��3���~۵��<��������A�]�p���"X� �g�� 6>�y�%���X��|���Vx����9{i�q�$o�Ic�
%<���8���� r�t����I�i6e{����@��)$�1�YH%cP�/��X���� �ݎ��\��7L��Hy\#��2`� ʲD<{\	��u�z��pP��x�t��L�Z�����/� ��~��P�y:x#T���w���#����T�5
_�P���r ���D�T� g��b��w0�1�o
��5� E�̽��	"9�.��חt}j q��,�������8B=�|���0���I ����;��Y��L�p��!H��肌	D'�n�s�Cڜ	Xԍ��`�d��v��hk! �� ��bXC��T��'`���m� ��S.(�v6	p�0��a9�_% �xD���g�������& �%�B�`�.О繘 FW"ۆ��,@ 
�Ñ2��S �.��ڧ��\��0�\^k+:a4X�r-���Z$���]H��dL�W�1��6/�E��^@�]��@�2�D� {�X��t`TC�*,v�� �웲h)`Xpq��%��=a�rU�!�������;���� �'��`��(���4�	�!�B�N��΀$����k�q�j����@� &��BM)�r W5+���}��� ��G ����]4�V�O����׫�?�v|� .�X��0x߰`����Y٣\a�0�!Ɓ ����q��p%w�� x_M��\�� Í��VU �D܏(`0�T��� ���K���C�	�!��� 9�x�����y���M�^�4m�~�SV�S��߇���q�x���oQ�P�m���ȭ��F �6�����#
�ߪ\��`�x`�2y�u�o΀�ˋG ���Iex�ǡ
D ���� �����L�X�8� ��W_#��������t�H\��A�x�q.��ߛ�+PU?xG7�^�&�����J�G�_\��z0��ê�@"v��f�I! �*v��:n ���C~S��w 51a *����KF�"����G�e�F�� m� �F(S��۫`Q��z;ю�Z�yU�1�{w�KG��P@�m�5� <.�}X_]��Mx���E��/Y_Ar��X ���נ}I�8K�ዓ��nڏ�~'A%͖ �v!)�/ �*s0I- ��$x����W�D*�4���("��Z���m��t=�#v�1H�+v}�=oP����U��0���HT� �u�	QZ� �v�HX� �"�d�� �[��?��9�Z��(�HS�vP �>ݎ�	/��X�HD�̇< �@�paV� ���g��W� ,�$�+��M���� ����0�d �mt��{s�4 �[�V^��-@���E���rz� ����\�Z�u�E�}��� ��VB�<�"�%�Qv� ��;�2 5�X�{�[� P���"�b�MO�R���s] ���쬷N�{�wȘ?�G��#���`�[^��H$��pL�� 8oa�{c�tG��,x�����Z����ɹXpDa2��X ��3�