MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �Ed�$x7�$x7�$x7987�$x7d7�$x7�$x7�$x7�$y7D$x79a7�$x7T=7�$x7e7�$x79E7�$x7Rich�$x7                        PE  L             �   @   �             P    @                      P    ��                                XQ  (                                                                                    P  X                          .text    @                          `.data    �   P   �                 @  �.rdata              �              @  �.rsrc       @      �              @  @                                                                                                                                                                                                                                                                                                                                                                                        UWVS��I��ŋ��   �\$�����f3ۋ�@<�PЃ��r4Y��	  ��APQh/o�X   TTj@�r0�r4$��XYX[^_]Q��U��`3��U�M;�u
���u�O��+���2B���s�5 ����ːu����А�D$a�� U����`d�0   �R�R��}�r0�   f��f�t���   �u�}�<Ar<Zw ���j �E�P�r���5��ju��B��@<�@xÍp�}��   �ë���u������B��j P�9���9Eu���U�������E��� �Ð�D$�a��                                                                                                                                                                                  S  (S  :S  FS  TS  eS  zS  �S  �S  �S  �S  �S  �S  T  T  .T  =T  JT  YT  qT  �T  �T  �T  �T  �T  �T  U  U  U  $U      9U  FU  [U  mU  �U  �U  �U  �U  �U  �U  �U  �U  V  V  V  &V  5V  ?V  QV  oV  �V  �V  �V  �V  �V  �V      �V  �V  W  W  'W  ?W  KW  ^W  mW  W  �W  �W  �W  �W  �W  �W  �W  X  (X  <X  LX  _X  pX  �X  �X  �X  �X      �Q           S   P  $R          .U  |P  �R          �V  �P                      S  (S  :S  FS  TS  eS  zS  �S  �S  �S  �S  �S  �S  T  T  .T  =T  JT  YT  qT  �T  �T  �T  �T  �T  �T  U  U  U  $U      9U  FU  [U  mU  �U  �U  �U  �U  �U  �U  �U  �U  V  V  V  &V  5V  ?V  QV  oV  �V  �V  �V  �V  �V  �V      �V  �V  W  W  'W  ?W  KW  ^W  mW  W  �W  �W  �W  �W  �W  �W  �W  X  (X  <X  LX  _X  pX  �X  �X  �X  �X      KERNEL32.DLL   BuildCommDCBAndTimeoutsA   DuplicateHandle   EraseTape   ExitProcess   GetBinaryTypeW   GetExitCodeProcess   GetLongPathNameW   GetModuleHandleA   GetNamedPipeInfo   GetPrivateProfileIntA   GetProcessHeap   GetStringTypeExW   GetTapeParameters   InterlockedIncrement   IsDebuggerPresent   LocalCompact   PulseEvent   ReadConsoleA   ReadDirectoryChangesW   RemoveDirectoryW   SetCommConfig   SetConsoleOutputCP   SetConsoleScreenBufferSize   SetEnvironmentVariableA   SetLocaleInfoW   SetThreadContext   Sleep   TlsGetValue   _hwrite   lstrcat USER32.DLL   CharUpperA   CreateDialogParamA   CreatePopupMenu   DdeSetQualityOfService   DrawFrame   EnableMenuItem   EndTask   EnumDisplayDevicesW   FindWindowExW   GetClassLongW   GetDlgItem   GetDlgItemTextW   GetMenu   GetParent   GetSysColor   IsCharUpperA   IsChild   IsDialogMessage   LookupIconIdFromDirectoryEx   OemToCharBuffA   PostMessageA   RedrawWindow   SetDlgItemTextW   SetMessageExtraInfo   ToAscii   WaitMessage GDI32.DLL   BitBlt   CloseMetaFile   CopyEnhMetaFileA   CreateDIBSection   CreateHalftonePalette   CreateICW   CreatePolygonRgn   EnumMetaFile   ExtCreateRegion   GetBoundsRect   GetGlyphOutline   GetGraphicsMode   GetICMProfileA   GetKerningPairsW   GetMetaFileA   GetObjectType   GetOutlineTextMetricsA   GetOutlineTextMetricsW   GetRasterizerCaps   SetColorSpace   SetDIBColorTable   SetMapperFlags   SetPolyFillMode   SetWindowExtEx   TextOutA   TextOutW   gdiPlaySpoolStream ��Ji}�����?,�mʘ�a�뱑��E���[��l4�����ņ�}���NI�W��̀<�`���M"��`�(#u��#t����r\��?���Ő)�+���"H���*`�    [��F>@ �M   �D$���   ���   3��                                   4&�kC   �vH7B     @�@d�5    d�%    ����g>@ �̐�   1�$�T$��1+$T$��W�����d�    ����㐹   ���g>@ �݃�>@ ��.��ѐ���f� t���؃���ܓ�>@ ���f� uܓ�>@ ���f� u���a�   �v��������Ĺ}�?�<�k/���d��v|lLDJ_hv���H��3�<�l�0����C;vة� ��0&�vک��}� �� ��76[��C������7fm�w7;��7/���6�R�fm����	???h��Z��S���<   ������   ��3����3�������@���+�ȋ��@JP���K�����u��?P᪯OA����@zO�?�@����?R�FiB����On����Oe@��?�)�?"�٫�O����o����?�OClX��OFq�E����?�'��[�E@�(�OF_�2ȯO��V@�F'OF@vOF��OF3��E@h49�E�2qa�)I���c�����)�Y�K���[i0�w�Ɓԉw�AR�{C�=}���Xt�L���i`�䇸�\�$�r��_0Y�XdT�.Jw�C+�"&u�е?�wW��'B{in_��θri[V{�����y�m*m��(�0l �B���?�`Ik
9��vv5+k�7�q% �hhAp����e\w0f�~�ZyK�xs������,���5D��HRa����G���@>�3%�����έY��) �2r6��v��Ϲ �d��ģZݣώ���ק�y���q&���Ɯ��`�]~d���%�1��NzJsx��k_��c�T���RD�0M�<��")�t�g�	�'&�ٹ	.�*O2�r �_��ty���8vZv�pq,�P��
���b1�C��r��!���	\�z3�$p������r�KÀg0��B��~Jo��`�V�W�O�/�'}��괒�z���I�D�d�h��p$s�p�W]��Io�(� l�Ǐ__7����Y6�MH��
{F�a����z�ۓ���7]+F5��q��2��/Y[�p�j�#��X���_"7Ji��V�"��(��+�vU����-�mF��pf�T�@�7�M�4�f	�q�Q6]�=�l�G�A�.�}��Sb��H�sۮ9I�D70j#�k�K$�B���zӀ�0*�M��3V1�T�b�rB���0�j��^!�>Q���D��Fo��Z"�Sz�Ǡ�������z9F<O�c����9�27}�{;NX|ZE��ˁ}�vly��F��w!4с	x�WO�h�L�o�:ţy������``�t�?�Y��T�zd|P,L�
GAU�죌~�E:i�,~�Z!�U?M�1���{�[��e/�p]��Мt݀u� zJ��:*����_`^�#�=	�ͽm(E�C��E�^�pmo��D��Gܻ�ρ�C�N�H�&
�����C��`�[��pù$�-����/}��v�8�#/F}��#�)���ģG�b
U��-���ݱ ��[=�.�mM��9b Ο�����rI�yR�>+�ѫ@2���W3�h; >!0��+�*x�����@Y��1��(�� ���mϪ��������n�%#��HSSp�1��@�Y�+~@�^j��I�Є�%����YL/�3�i�$�q�T>�G<ÄǪK2U�R�t�IdAj�[�eL
aF���
	˫J��@��BN��S�'�8l�,��UGk� ?�tQ���>.�׶�G'-�^M�:a>������ݍ�����$NH���{�V#�H&�$'mTC���լvZ�����k�I��*��E:J�1�R�t��Q�CҜ��-f�e�Tƅ�--�b`#����B)e��w�6��mI�5�)i���zAXy]E�+�ݗf�ʅwY�%aiS�R��A�'�l�[6t(���c�|'ѥ�kا��s&�7P���U��p��{������l�9a�R��	�"�9����T�[�pΆ�$2�{+��v��QmZ|COhU�P��q�n��C=m���9,WCO��l�jm�ryV��k�z�,��ы����#���������3��
����)���a�Y}�8\Q��5g4�sH�v�'�q|!g�9�M�@���R��Ò���1�r�hF��Rq�*7� �'b,1��&����o���!����j1�o&KME�?x�K˕v3-A�M����s_��v�\�:��,�nA����\&[���.½Of����T?嶍%e)/ps@$c&x��*�d�Ճ0{���=�y֋�}\�.fT}�����SϿ/I�XO�ۯ~*�n�Z�p�:Z3��!�N?���<4�rd��	Z%�C�e�O�vz�J�T�<��m���ɆB����G!&xۈ�Б_\.�a�f��OL��A�!j\�+�n���������Z�^�1`���ޓ�%��SO�aq�6s{8��hqt� ���e��MJm�V�^lP�xh��y��;��#&�k�E'*D�%g.k�u�ak�w�}�~F�ýd���hM��m�}1Q�۪�{��o��ͅ�+{!j��-X������#����K�%y11YN�o��c{K4�˟�Abl��GwN^0���4��X���^z&��������.���YAGjZ:alxi�POM��>,O�٩b�����MĐ�t($<S�w�LD��~�^�2�!(��IG�+����}oK�S�uqI�5
X�#���FB��< ��K�q:���ڔ�4��������W`��[��3�����id�u���Z�Į���m5:W�R2�΀���|�$v"j�֪0�m���g#�A�hyt(�v�ɪ�����l�l����y���^r9Kc�7$�fZ�cg^�_�:W&JѰk V(���>]��4�d�%�u�k�́f��qޭ���r-�+H��W�.�	*+�E�v.���L�+�/	UEwj�!f%V�]��k��(�L=���	��C��0�+�<(��aI��x�rpR�=�����Z2K��V���c� �#W^O����4�8���3cnUO�����^��?<��:�-���^�NW�QÑ*�ɇ)(�$Oۇ-�dn�r@cqɞ�3h�������J׼n��W|B�� W�bt;ˣ�rK�����?F����q4��i�,�����{��I��
�����2�N-�UG��X"X�|�+_EA�-�N{��,^���7H�
�ȃ�\������
ø3:�3�LL�q�L.1��jQJ]d��Eˣ�3��u��.��4��7����b� ��p�dl ��(��Z�-�Zo���C��F�;x͌]�'�̗�*Zh�s�\�4QO�������W�1y4�4�Q�����'��hf���H�#Ǳ1�ʧ��W�F�\��M����m��P��㿈]�M^5a�=6�J���Rm�2���L!�m�����mݷ�z�ߠg�GAN�%�vW����Ն�O s���7�bDL�!N����P�a�~���?D��Z�ec*7�L�\=�5���֤��/��g�L��!�y�u�X�/L���Ġ�u���U���Pb֋���1���>]�k�9,e4t��,)��ˮ9�b˷���t/��]* "�`����(֧D?�Ԗ�+͒W�"n��D�G]�Ù|�ޯ[��\���5�΢k���7 �x���Q������qp~s���ل#��R��r.x�em�L�x"F�+�E9k�2��u�~=X�DH7�T�6R���|�^��s�V3!�U�zשj]������1�_=��Y�4��u�kki���I���p@��)j|C��{�7�B6{�f|�I����G�<�e��{�tS��W|MBU���ş�Я4�u��u��ll㇯e��M-�A����1W���b�[Ǒ4�wGn���7N���f(���}Z&�"������	�������FKhݢ���EҦ�NRM�����̓�]J��n��s����B
1+�����\�nc	��/�d3���$;��
�V��Q�i
ZL!w&5^�3��%��}����-�ޕ�G�][y�]�{G�c#��F��S%-��I�*�.%x[�q�t�"d����
5��,[�L��$X�����(��B���� �Cđ��n����҂ڔƏU�t|G/^�ﻏ鞆de D@���wb�����Lb��� ,�iYC�E3\_��_�t��\���A�b{`������w�,lU&���^���>��&r[�8�z���y���)E�{�
��mb�N�*v����Ä�Rv�uJʻ@D�8lt��]Ey�v��Q[��x  �O�?ޜ��L�I's��]�
���ѽ����C���[u��z�n��e�k�j,������`c����1���j������$��a�n�<'H5�\mj�-���<�3�� TE.0SV�	?.+��w1�F]�l� ���P��l��Ѐ�q�Q/]��uװu���|k�D�c�c K���FӸT�,��WRC%_�7N����2����^��M��~��p4��T�ள�v�3���V.`����[�+(���@��ꎛD(��r�����OJ2��bZ���ad�� 4b <�4���ƑKֆi]+M�*1���ADi����>�q
f�= t�lr�ܷ��%�S[���&�Y�@J��e��+rXe��6�㥥�%�7h�]Y��Cy�����*�5�;v �8[(敢�ωl���t>�Zs�^5EP��[�ߘ�\�	��(s�~�yZ�[��kB�� !�t��p���X簨"��/iq��Mf������K0�E�f;αd���2�0 Eӌ�Ӻ�=��}A�&4��^?�l �����=�k�g�ӓ���U�g bI�i^��p+��ٸ�8ͺ5*Mq��r���0���K��g��zݗ� ~�$xj�ד\E1�p�>�Wn��X��!MPt�iQ̝}��vT]O�s���:�Q��9E��)h�`���da5q���"���,�o9o`,Р*D7�8,��z�d��^��� �kI��[�`�< "���98�� �UD�'jayZS�vWxV�Yj�� ����d�(�VLU�i<,�#[��[�̨XOT&��o��!�bB�?�oO�3%���o�Je�.�&E�9��HO�m���}B�ʄ�)�6��P���27�D�K�q���Nk�o����8�X��힊�ƻ����>���p�w�5��gp밫�aМd�{�<z�����qt�KT��W�ӻA\Х+�Z����/����� j��
�1���h�3,��:���&Fu^��/r��R��C��;���t��T�:(D�
�C�@�LYgͰ����?�r׭�IyɉeN%f���S�"�n�����Ht�������p+ݿ���J�������u�Lt�*7����y�2��%�m#~钹G��fr-�B��6|
���8K��6:�ڜ:Љ/���W�;�����M,�_<����'��V�M�׫0.�l�_���ty��ݤ}8��jA5q5�sU[[3����.=h������~G����;Tf��a"^�	Bp{r'�4%��ѱ���j:��0.Յ#�~��l����b7�Mk�᭞���-�XK�֭�k�'�,�b�}�oF���]�0�DuL4�S�smx���^odI� �:��^���� �w>o�oG"���43�z"��0�|��M0 h�.Ro�lϝ�P�-�=��y���˝�"��7G�!⣶�J���3N�K�1W����Y%x�8���C	��<�/V�E���a۬���֓��U]t�;��c��k��`��·f��'R�� �2�ò�͗8d�#@>|W�,�q9j3Z�N���+-p�R;��E�؜�R���'�K�48���T��R;[�O�%���Di`��ZŪ\���0�^�ۢ<���|i�*��*�C�!��4\�G��mk�+�T;yP�m��1�oտ�1;#=���C�P�G���Ê5U$���f/𖖦��򯫧��@�ձ(�Y��J>!�������JId-�ՈC0Fl������9��9J6��1L?�Q�w�]�}���tگ%ٸT�O�ׄ�.D�X��P!=v��p�BPpR�"λ�T(T���,��۪�.�u�U���v�P�h�߱�!$b�H�=`�np��^�=�o� ��)>[z���L��Q"{�h��o�a4jA؛����1����� ���*$t��Qq� P"z�R[
٨���.V-%Qɘ������i'��4̴H�6v1��s��`5�.m˯�5qE/��U!y�� ee���"�KFFI�U���������J�h��wHy�S#��{rZ�D��0���
���ߌ沈&������9Zj)���.a���ȭ�w=��t ���D�ì�O�d�%~3���I�\<s/���f�¯�[0T�������|K�N_Ù�� �_����ԃr���qCc�^�y`0R�F��0�p���vL}q�8|������q�����6�1����i�Z�f9��9��ܒd�7��>�Zc�$M�3�&!G~���~��"ԶDWҚ�֛��+:��U�`#���w]_�-�P�n���]��.���]�ǰKƚ	��$Q[��8HK|̈Ut�3�H�� ��Ѳ�u�f ������ſٜl+��Bm$�gv�3��Eȅ������]�#e����q?���蛵$!Y����?�Q? �t��n��c������<�.h�~_������7�HYֳ�!Շ�4.%u�*���3������᩾!�k�����v��t�d�^��������,7� ��4��?�e�w:��H;���X�4��!�b;�M�#���R��"�3�\yg�𛉟s�����N+xo<�F:�WW����>�%���-z�������w�ȡ�yt��F?<�Y;�Ú�,-�L8WI�C�R��*�T����j�tp���[�%b��C�	�6��S�Ŧ��]]�QV��ᧈxJ��-�֘*B1Tf
�ziAd@z`�J1��I�K�t�!qD-�)��V���#�>:ީ ����o�����}ς��"�8xq�3H���	Z.0JL]3R�s���
s����>��>T	�����6"�DX\6�m�@�o�<�:�?6J��yvp
���0N��"}�q��)V�M�aA{����UWG���Op3�j����ip�[��$�'JU.��9]��])��3��1���"��O|��=�<�W����#gQ����[!U�t s��eO!�'@W�F�3�m��K�D�ºq��e�Tc:�e���3C6n� =t*+c*�9
���p��{Ҕab�6��u¸�C�I-��j�m4	}ʷ>�Ī"��)y�R`��^�39C>�����r���ʙ�'�KSK�����F���e�wċ�"@~0r�r;暸�c5ϳv�W���t�6x�R��i\�r�V�� =�HlB@`;]�7>:Y�F+�tw�ο����)ܰ_-��]IW%�{\�I����kW�B+�O��;��%�rn���M��h��k���`��𙳂��=-ҊRH�?W���U����>j^.P�S4�g�niMP}��`�{v#ȶI�s��sdl�u,�H����|or��C H֪�9��&7d�.��!^�_ �Õ��M�s�G��Q�w䯓���f�@4�,68��	oz��`8���FZg�Y�:�\8�̯��u@"�к�%�d�������+�9�(�5Ce�p:�Bk	�������	ֹ{>?-h�+"�Q��Uó�g�O4�ܤ'
p1�ɖ��u,hO�5:'mz�Sta�7!y�w��XB�$$ypP�e�si`�0+�	�s���i����p��\3�O�#�����z����1.}��B��9����~ᯂy0e%{k�!6`��D2c�����6@�\�P7�1��%"q$ޗ.2��	_��P���u���2���1�!���z������4��������(�ϫEޝ0�aO���U��r�:1a��3��@Y�S�9u
�B�2@Q>h~e�KB]��
�.�~�*������������v��P�\��us��N��/���]#���=d3���_S�k��k�r�����:�00Z�笋��֍JI�  �d�kL�m�b\z[����3��c^���&���2���X���1�����i�� ��c��$�g^���s{q��6j_iI�tct�xH����4��B/��p��m��&�J6j��c�F�ߙN�I@B�������(��jX���:��p�h8e�GM\�ۨ�P�z�/2Mn/��G�Z�������G�ׅ�˾���	�~��ut�wƮA$�o]�Wj��l���r���U�����[��T�}M�d"����Q��){5�^��G��J�9"e�-�w�D��+��y�Kڱh����3U�!R��G�ώn�K���h�<��\&��c!�++ �5f���i)�6K�^��z��؄�xn� {~q�.)���r��}L;��p�rE1������t����)@#�탰=w�|CLg{�.�X���~.�+B-�6!���^$A	��;��r�MV$=��8Oh�t�:v��M�h5 cc�"��~`�c�k���G*�?ܞE:����8�J#W	�Pk���f����X����Oz3H��n?c���
�-���FJd�j�{�v�| �ڙz��1�sVƋz�,�������$t��� ̮�6�������ǵ���!R�,�t�C�7<�H�-�8<	�/�'��>#e�Z1W��Q~c�L��yHs&ѣ���"IV%��|\��D>���ي9��V\v��>8Q�@O�������%ͧx*Z1-��p.g�m<�f}��JQ
�O�B�R����?�N�!�h�\&,5��rBW�{v!�a����G�v�!��.�l~�R�'�����wӲ<��k�\躕/	�9����}��s����!����73jr�T� ��W��r$���,�{�,~�#ا��S��{QuwNƐ��Z�NDz�Đ>�%�����!����^ϕ���J���?����f�rA3c�7���SB����}��m��u6��{�^͞��Nu֒苙M�>�Q�[���K�t���d��7R�]�������O�*�V�aN(;αF�ά	 ��;Hmalm�c���;��N�v��|V/�[���P��G�}geq����?>��dj��vn~�U�7��2�$(}�F��^�_̟O�R#�t�YQ����w�n��!4&j��^�H�!ti����tnGx}�yx�j'��T�=��+Sm��=|�B�O��/#B����<*�����,�b�����FS�Q��\QGs[F����d��礖�����.M��t>�W�(�3QrhY~��}��禔{��T��E��ɯ�ꮚd���8��Oq�ͺ��`?�]F��[vonh��P� ~�3�Y^.X;�S�&�8h�J��Q��(�	��I=�}7�/�nWO�SY%VNZ(O�������,������~���$�û��͎�t�B�@<�VX%%Tc\¸��-XLC¶Y���
Xr$@���*p~�܊���h�V��S���/�N|Ɗu�Jӟ̠M7�:*aG�g�u��zޣJч�I��M�#�ϸ�B�b��Fr�p�@��<�M��t1)���7'�-�fI���5�M/�j:��DK�q���^T⏾���Dm�<g��s��X��b � ��!��};���\0m�W<��h��Q����8|�D�K��'���=Ă_i�J�K�U�VX�jH���� �K����1X�����O(ia���,��v�|x2�Ió�����MB���`'V����5ϸ����*O�ĵ��M�`D��d�����q��6O���4��)��*M��$�؛oK0Y�9�ɡ��rǧ���2�Q��A�_kG�r� �������!�PW�v� �H���J�I���T��S�c�@�g�,�- �WB���5?���`������;EKh�e�,��R� �r��$1;S���J25+�}�]E�WA1�ݙG�'�K�PF̒���/T�����&�R�/u�YR�gO�=��?������-^�e�1����e~	�J�_�+�h.�E]Y��W�^��8؍*^�/�Nx��bld��n<��QAHm�d�Ιm>�[1J^�`"W;P��nA]�����ʁ���F�6*�4X���f��4��:��L�ߩ%k��H�/�N<Z��lʨH���xKN�Cْ&���
���}n��ﾏ��Aբh��ͥ�z�L�8����u��[о��'Jɵ��b�t�?��ҵ��2��a'�zZ�{�SK���9������i۠v��E	Y	6�x疘���-�v��E�i�b�xR�B�
;��aB��e]�]TA�D�1�\�%E�MՖDQN�O����otkG���U<X�\�U�P��#S�qq�OD��̾>D)E���V�Jx���[�Y�����I�g9���Ii���9b�|�����8�e,s�"E��nN���-p�̘�T�&-�(�Y�	`�]R���B��O��=8{��Ois9�{�2	Ͳ6�@��ɶ���h�yL̰K=�
�U���U9J13UziUh��9�㮄�*unj�� w�<�jϖ�NB�>��}�_i�����v=Lh��y�bE���P�q=�ƎT�|�;�康�^��o:���5D�e�_d�4�z�J};3R]���Zs%ӻ��bU����K����~�	��ch��-"�iڲ8�zX�?�)��.����t�������e����e`�sg;ϑ0��˶�P
 Ƅ�@٬�4�Krv8U��D�mb�W����8x�r��S� �\�b919�]8��f��K-�[��`:Fק%J�^�ݰA�S4EAK�^��S����`h���ly0h ���zV��0Mj��C��B4b"Ɓ�4t+��9fΊ�x�1?A
�Q�b�ZY��Q��9���wN��V�ț��~��O��"HhXZ|d��m1�MȈ
<i4��5����w���d��� r%� G+UT���B�s�{_�]�O��z�K����#�+��2���T��3X��MU����	������ى�<[��5*d3D�T7�[%Mݫ,N������C�p1 �':�z��S�Zjo��"^���Fm�������X��)͠*��n�a�e�M�\��:�	�$]���Ӄ�PJR:��L�
L�$^�f<t��*r�̎@�-~�2 Π�Ǡ�Yq�nQ�7���t�:8�WZ���	�m9u��|���7?���C��+�x���ڎ������̃Q5�o����sJ��h����m%K���bA���E����Q*���$��:�I'�M'ҹ�T�Cob:�l
��*�"m����fx�=�����1��C���������(s��1���	�V�"桨�#)Æ�ŗg�v<fH絍�pNc��������O�l@�g/����V���[D^ߒ���5	�l���O�B�>}��`��Z6�*.��8�E�nEt ��6�b�&��x��ҏ��<��D��*��Cn�I�l$�f��OJ��ZG@�z�'O�ud�Y�^mA��S,�(�wD����'(�8�/�
R�<����<�Y5P&e���q��;�8��N:�����
Y�A=�x�c���](�1/��W*3��[�@���9P���#�;�!Dl��c	u$Њ�2�$^��:Q��DK=��jHS�~wyW~-MXD$$'L����� |`����Zru��-,D���RQھ.���xWe�u~!y¨���֑�2�f,�(`���x����A�YySw��U�4�+����$>�?Y븿��ۀ��tB��P$�ILX��� <`���"�δ��50K����k=ba�P-�Q���_�<��ջQ�;�lm�,{��!4 �n�h���ʙ��,7������`�Py�(��X�Y(Pz��3��ޙ�<�(:�`�&��Diݼ�P�Yxԩ�eֿ�/�nE-jjԻ�#^��+	O���U��:��yS�h�~�2�?P��s5�a��r��K@7�F��t����I��O�n\��[��L_���-���t �.B�#��G�d��BZ���,�X&I?�dlZ��Ct{7���ǺNRڇ
O��g��Íc.U�Z��!7�k�;R�
��Ppw'��X(��кv�&�~�mf[�Վ�EM����N;X�:��(��8t����Z
��4�d�v�����z=z@��}�-)��@|���9E�����N��5�Ka𹢺�tt9 ��D��ᘒ9�eЕ3톱�U�S\�����F���-�a��l�.xrf�0|v߸��f�s�h����s���`ɎK{?�K� g��V;��+�U��ǟeC�d�u0&A�Ǳ{y\u'�ϧ�&k,��5'�S~��lE��kZ�g4C�;��.�s|���v�]��^�������E���HkW�M�������@�AP��@1�P#��pZL�sr �ع��PF-��d�ċṿ���mn귈o��T�I�%��\�-�X�\h �L^�XY��C1Lw@
�A�+V85����5�,�so�U7���#����(��tQ��:j!X�Z����P���n��n����,U���5��I��f��.Ѐ���;{��5�vf���kZ�%�c�ѳ����v���N�d��7\�|��ڞX>ݻq�M�"'����ž��xt�"*�W;����v*��-G�9G	���r��^/����p5NtRq��U�A~diVD�#:Sm���&�-3�wVU���^���r%*(�&6�~���]�M�X�a?��ڞt��Ȇ ����a�^��VʊKT�A���@a�Yl9��~o�.�b�H��=�����=4cL�s���;�ȫreX�4��"W�J@	�d
�c���"�R�R\�̜d>(A���7�ŗbN-5T�]�x�B�Șߋ��L���nu|~c�R�l>�o�f����/pޘCu��Mp�.�}���gQ���H(Wc����[�~Ir��k��'�	�����.%;g�:P��9���Y��5�dZFS0	cQu��u�"��sj�R��� ��0���+��n�dRy{��]ϋq�|�q<n�!�*��wd�M�t�J�f�o��a�{�>���F<3`�1Y���O�#��"3����D�'���[��-�zĒ|�7��'p%  ��E�(�S��9��s�Ή�yx8Gj�\+�fؘ��S�=��C�G���|@ nVH�w��w�K�(���F��m��!i�S��5��L�:։���Xp*����=�w3^Q�Q�/�|�?�$� כ8@J��_���cQ�l�~���X�s�e�F�5���mT2L7��s�^�n=  Δ	����TQ�/��O��,ۨ���vd���2�_��Ҳ�^��t�gO�A��e���jS�'�������7y��gh�J2��ze�)#��H	��B��;݂ړ��`�w:2." !x�=�Ȏ;�ӯ�W��ڽ�ՄqU>"���]�T�E7T��L�Td�R���P��:@�{ĺ������X]sL���)�I(B
Aa)�|��� �70Ǟ/7g�%���i��>i���%���ٯ���XZٙ��X%�	�S�D}����8���n؇�e���0�� !떴��!�΄��##������]�0��`�E	���/L�5;5�i�0m4M'�MJX��un�pI��t����3
W')B���6�R=��u�5G!v]"�:�H�"������6D��NGi�&��v��RcHW:���ϰ�ғǅ/����6����U�QC���d�Z1���Q��q4<�4g��Ο�ff��,�R�RI_�� +	O��qخۓ�7�\���M���H��f�Ȱ7�r�V�Ũ(�r���?�Q�c�+j q��X����B����<��9Ч"��q�wE��`���pý1��
V.Y�sG�9<��K�������Yp�$���Z���ٙC�}��x�ݴHC��H�Im�~Z��[ھ��%����]~[H`�������%Лa����NK2����U�,��k"P��y��!�W��% �r�y/��&��J^T��c�g'��z�s�;Zʪ����:j�Y4Z�l�_�$��:�A��a�hUைG14�\�Ԭ2�2�DHS�����i$����¨c4�� srfK�Hl�pv��b�͟��\�����+k}5�f�X}�[�_��'��i٢��mH�u���{�3[���kAa�V) ��p��yH�,#,�)��n}v��7b6;������J{���\Y(�/�z������"˫$�z��V2v��]���iԙl���L���j��[�	1@-ujmg� 1��o
C�"֢]��%�R���n&��7�?�e�7�j?\�8և��/,D 1.��ѝ8�����~��Bg���Я�B�򸽌�5��g�(|�I6�5i�o7����qn�n�8��Xi�Ʋ���`���F��u�XT�W�.�N��2%�);cc�Ԍ0�g�Ǽ�����
�(�^��V�$����mS���z�$���!�qb�1#�;�[���&�D��nL3p�#�Q�����<U� ̺��~�^s<BI(�u�jK��E�4i5������P��@��]I8��V	�C67 �Y����xhzy��ہ\B.�3*5Z�?~�5�W�T�5������4���5��A���V�(�~ܨj�T��}�<#�RAR\$�<�Z�#��I5W�����J^�kC�8wQKV���*��Jc�MW�rߡ���µy�N'l62��B�CB�E�O��#X�WU�# j��qǁ��q(ht� ��%O��8 G����1|����#���ۯF��}�4��n��q�ب��F�[�/E���)����Q/��$��'�M��"����\#���5�����T8
��<���u�"���ljgW��]�n�0�䇺�3}�'z�^�R#%�p��m��tg������%D%����I�lA��j�"mK��,��`^�J��q-~���@ L�c4$`�	�T;���N㶇-���Hi`7�@�]P��U����^�Yk�g����bl�~�D�&��s�\FT-�ෙV\K�#y�j�/jA�yA��7�	�P�r T����-��$��{t�e�F�N����bn�Mh>�W�Jms��3���R:��T`	����%���-PY���'�D��(�a���������`����p|�
�!�g����i���T=�����gX&�Λ�&�>������3�Z$l�6T��.Fr�6#:�l_	F�Y�0(��-�����b�������`8�Я3P��c:�<0@��4��v'q�so��iX��ִ2�ys�\�.d��[��n眓�� �<QR؀��b[�;�_r�l1�zw���lq�i5�i������ ���|/A+����DW�b�'J�e�~F�@ɛW&u��_�b�S���-�Y�h�����-R�0L�Ƚ�j��Xi����/x�c�8�e��i�3����J�-R̦b5l�ރ;�X^�J嘂J	�D5pw�D�w����S��4���wmvbA�~�bp\�����Aq�o�q�0(@؃v�@#^�.:*��xMC6�� O�����W^������#ϕ��������Sg�����zt���^m�嵬L`"1�w�X�S�%o���b?0B��c�#��vX1�/w;+P	��OL�щx{ ��5-�I$��.���H��>��v�*��� W�l���f�w��Xl�]�J�� ��� �*⺗d�X5�Q��4��08 :�tF�z���r�A���T�5<�w��a0�Gȧ��_��� i]M\����0ػh�c�O(��W���$מT�c)p}����+�X^4�S�ks1�`@ޟc��Zz5!]���YN��f�7��1�p���Ys�d�i�O+�Sf���3�%t�Q`�����Q-U����ռK�2]�7���O����K�Et�.�I>��yxn�(?�.��0w�K��Q��H� �g:�MrȌ�1�����Fg����+ާ�9��<�z6y��n��F��'b���ӿ\]/�
P��7�y��0\|�d{f���QED뷿?YZ:r���Ξ�3�S�`��,M�>���c(��%7�d�~?�7�vGf\��}3�+�)�Z)O��\=�w��0��J	�˿w&+W���S�����_G��D�#j͛�w���]l��	;E�b��@q6[t�W6ݦ�����L08��tR����#���-4i��>G�������V�E��6�0��:_�����aE/d�7NT����P� e=�ka;{T��/C%/F�l��]Ub��1��jxD�� ӠA���B���|a�{-I�?
C�t�p�
�{���1�E���"x$P����:�ל&f�߸*�\������b9ވ��x�����O��&����9���Z�Z"�Ҏx��G�cԸ�ѭ���^#�a��u��ƲH�p�����X���sd3�]X/��{�[b2�j+azQ�`%LL��)���8ȿ,��([�_�n-�M��\>���'*<��"�N�ې�C�uy��6�y=�DY2�`�z�x.����ͯ[|bܙ�@��Q����[j�0K��iH�Э Q���t�JZ��C�NM���*�i��&� ԑ.(��ۦ�N�ű���{z�.�����þ.��	�����s�Q�ðQ>�|��ZI4_����L+>�����{��-�&k�y�;�b&�����4�ʏӁ郃5P^�9=���cQ���_@,��2|���_ד�A�#��'�� 2��${�������¦y-K����ؔM(�|bh�����pйz���wd�y����ɍJ%J(NA����W������g���������k\���ݨ��O����o�����t������i�W/f۞�+)9��YR�;�����Ѣ�]�A���p�]�Ӻt�+�*m�F<����k�eYܭ<#[�r,�!�� ���ϭ6hO������`��!�B�:�!b���;�t�Od ��:e�v�nɏV2�
Es�~ȧ�I���RRp��0A�Y��r8�e0[v[ ��IS���X �6ՙϩ��a|y���L$���Ea�V7-k�ցg�,����-N�������f�#0����� ��W�I�e�Z�aQU0�梁Z�8��2�m�/�n�\Pb�I���]K�Ua��z��7���~(�����%���ҕ&�h�\m�h\x��@��	�M:'���Qg�c��S��Z>'C��c�$:U���H�B��� ���o��4�!ï��<9������C��'���8+n��R�I0.�hݚc�:VXBZB<�!L�b��*�1�\��'��S^'���/�ɳ�`ďK�^��a� ��ӱ��N�cF3���"`����g��T�~٪�G2���7��.�T��E�K�j�oS��g���6���)_�6��?G�0ck�\/���x
VH�,-�!�O,����jp��Z-+EU�_���ijZ@���[����&h�9��0%Ԝ�L5d��6�ý��e*�02S�"a�m��G}�$�/�/h��U�p�D�]�/E���N�Aow��J�䆰^6\����e�O�K�p��������]܆��_G9�M�����b�Ia3,���{��PF�^1W�e<�s��dv(4�H9��(G��vt���o�$T����:�6�_��B���y�]&ͨ�؃��䂖�03Ry2gH+�t��o�� �4f��_�K	L/y��dN�hw/�C�#�1�7[�?�ai�J�X�O��@89��&�.�cEK�V�t�Wh����EZ���+�6������g�ߩނ��	&~���~��y�' ����s�b�U��ѬE�(�'|��V�N�8��P���+�%����@9���BZ���>E3L�ދ�&�bI���vSV�(�t<��w�S�/��v� ��M�Qk�g�S�z'5�o$��Ik)�i�����eTܝuv�|� �`�r��#V"h�X��Zu���ÛNUJ���	,#��n̝���	����I�!޹��O08�Xl����M	=�z�`V��1#�2�(J��j��h&i53�?�s=J�Ns^:��_�0O�����X�`,����s׭����C��=݋R�4��m�%���8u�D�Ʌ��&b¤ř{|[{1®r��I�^�1�	�(�o��:[� [b.��t���os��5�%)R�Ѐ�KE+�r�C��s�+���\��.�(�u��x �^��4���4(.����x�0v�Gb�G
pa�)�Ø��'���+W_�꒹��w'��W�xc�S;�twg����#�)�f1���͡�g�?D�<�����_Z� �G�$�<tU5t�8%0mw�(���Y�r��A��������@w.в��O�|^�'�Y[�`���zɤ�q�i-��?Yu4�ۦ��Y��?N�F�}��k�y
л��4�s踙�n�Ÿ	�pY��1!(�-�c�MzI���2EE�(��[��݉w�h]&Z���J·}�lN��!+��3į�J���м�}^�[C�B�߳}�eR��T�u*j �-Э���sh�@��P��xI�:�Ajj���H�@J��4��Q���b�	y g���#� ��WmmA���N0� ~.�37�9� P+w��h-�@�uu�{��z�:����%�*���e�
M�-8x�&�m��X]7���Cc9�V Kof:=���Rٹ�a�#ogPc#�f���͔gIL4iB9��>Of�Q5��S��r��g�-�~���^�t?8�3.��I�6x6�?+�[K;c��^����K?�=�;B�f����Ov�۬`�pPYn�������As:9	�JB��Q��	".��&)�(u����Ys�"�I����"�̞���aց!���&��9�|Kp��Q������\a>�I��d�v�7V��,���J¿0s�?8%��
l_'�~ż�)^��|\Tm�-(��$�$1K|�He �T�Tt�Щ �VBk?I����k�1�59���#����w�>�4+� ��5o;̪l�Mu�����u��H]5P�U���a�5,��� ��4���:ɸ"c^���a�zK�<���CH����|�n�[V�^]��uy?��?�k�9cDf���Z��?;�C�&@td�oUd����`Ȉ�jk�=�C"�M��Ap���P%5���ܓ��;�2�z�Y�dY��.��۶���;��0VJb�ią�H�a�o���%�mYj%b����.у�V��ÃR�r�&	H)s�]��uWFU8��r��J9+�oF���%�"�� �J�8��L����iI����zI���D�p�D��{�M�?%�7e��J�s�e�LJlN{J����`�����#�/�v�n|	 U�G�T��|���g�\J�����IT�Ӳ�zwJ�8�t��f��B
mIjz��Ri<��Z����N_s:�7[��6�^6階�޽&��hS���^a��o\=��a֒��^�IN⎊S$��]�Z�wTD�����QNi	��J�{�m�2gގ�H�s�<\��J7Lm��Y�B�0�Rǋ�v�*�싼����lF_2S0,�o8�m����z��F^�R��.Sʰ��	O��Qxa9T0� �$��)�D�t�B�S]������*����N��|8#:p�"m�F%��:�I��F��C&�[zV�I>�7\�h���0��Q���j�)��H]��߄���;`������n�����RxH�����P_��9n��.H�e��֟�ke�mt��"�~�ޝ�(�nJ�K����H���.jF[*�q��~�`C��	�ԘI(�½��xʍ���,Q���Ig *##n�:~��$[��j������}�c
Ө�7�����W���1�4+ܿ�2�N_���{12����I	��+=�$���)�֕��6Q�J>a��Xf����L!U%:P��U�۱��S+>*�E����k�N�����
C���	\_g� `v�td�f���arՂ?��\�/F��4�"��K�������m�>�Bx� �'2���n�0���,��"����"�2G�d���RT�oNI�3��_�Gke��{;���;�K?�<��.�,�J�g�W`�� ƚ��%,rGo���-ȾT����k�X%�*�|s���X_�nJ��&��We�J�ft��@~�O#���@��]\7I_�ϭ�ɟ"th���H5Å��V���W�Z�d0�)�r��фÊ� ^&�S���mrL4N�����"B�e���p~�/���i,��<f��g��Q����bm�m�J���q�&�G8/�(�'����]-7KG�\��</��` �&�Pe@<�h��P۱N�̱>�t�v<����M����J]�������T�DEؘ�����H���[S��%��A��0�����ʆ�ި�����=�̕�9��i�8&�k��YJ, �v��f��Q���0��[���j��C�6���+�0�f����;.2<�� ��&ܟH�@9^� 'q��ކ��u�QvI�Hu���1�!�U�����ԫ����YJ�F�FX�����y���[qD"@�h�����^�^��b�c���i8ᄗ!��qb�Ly�
�z��W
:���M��SqN qZ��%
���;
�J~ChdwVd��I�=��\Vr
�ֳ��e�q���ˌ kˇ���7˂����(j;�
�3�>�� 9.�Jr:�P�)`��S9�"�w�J2��V!�Ne�L���uO%1D⹝h2X0?3���\�wl�6回���>`����'-�����c�(q$Q�(p��#���N��I)���3ޥ �`KˤԿ���Z0�FD^ٞQ:|>�(MQ��q�w�u��y]��?S�����ڸ�7�Gf� �5L;�J|~�>�v�Լ�"T����g2XO���;;A��������f�N�=���{Q��j�=�`Z5�}�|/�6Ў�1��%m$CԚ��c(Bn��x����qZ�%�aJ�xf��1 Rv,QSfj$C,E��Y'�he�q�5&�ֵ*H{�-��z�u?[j��]3�~|���9}ſ�^��쥚�t�?�D[UPp��HN�ij3��l�E�X�Hp�a���WRn�uO4�f�(�?ƒ�_���?l�y[���g]*����fC+]Y�A���z,#��r��2�]�1�Q�N����>�"/��!��5CP3 �3������>��G|T,�����)m�E���#T%W�w񩞋��Ɲ��j�"��y*.��E�V�-����Us.�9ڜ�x����8����f�ڨi��p!���y=���k�ŀ R�:�v�b�������mt���%ʝ������
w޷ؤu�ƌb`���[�GI��ȓ�N�b�y��Nq���CY�^%��.j����{�Ǒ[	|,r]d��������L�Ɔ�^��#���f��-O�k�1��
V�ф���9a)_���#�@�L��p!`�r_S�ޢ
j��lw�i�"�q���O1Ad���QTW_�O��Q=�Mf%L�e��[�N��	w�⫒m~�`!D�Y7���$�s�Q�o����h�75�7�)�����C�F�p߯»<ǔ��ފ���d� �;���b��
���?%^�����%��mڿ���)��r�o��/�b�7b��/����ٔ��s�m>s��q�1{����ΌZ�ѱ^��9@q?;��~
�GhJ�=1Ԟ�;3-A]�k�|�r��E��YE�$���5�CF4�~���U:�N��v����Ȃ\��Ḫ\1ԋ^rv�չ��8^��M��|@��d�� 2h�H�����!6|��m�:��Ҷ��
��C#Y�7���K�S��U�ȃ��S${^30��(�ت���\䥮���M-V<��I��?!҈��EdL�s#gƨJ�v6�r-���8b3è�%�W�5���kg��� ՟�Gp�����ɚLB�n�!|�m}5X�3���:�iLn����?VRS�~<?�=���Аsq�J�oG�b�ʆ	��"��ܑz�*V�{���k{^�<�:�3c_؀��|I�%`����h�_kF���Ţ�]C�B̀���ƵE�� I0�I���W�d|,}��t��ò%��%��|�Pp����!�u;xN\G2�38))$��ʺa�z��&�j���B��!U�㜓F�Pc�]MJÓ��ƛ�.Q^A�x��I)�%q��9T���C��ٙv�����g8[54�#�k"Wegr4?�^����|E}��3���V�m�b��r��A��e�Q��dQ�oAL,��-~��X;pW�xe�r4�^Q���H��s1�:IǢE��V��ꆸ?h_.?��	�rh�I 	i��4�9��/.m�U�,���|\/�q�V�$'YW�Bӭ�n�b�Pfx���t�������D�ùz�WV�oC-L�{��-�%�#Z�&�x'}	'�L���N1ĢgaT��`&2�33����Q�u:��V�dE����
(n����՞k�=m�*��7���NG�>�z�9�6�I�#�U`7Y�Ǌ ��ϵ|	GrC{N*��be�ߥF6�9_M�%���� @��Le�/Q�o���U-��c޵���禀Q|4D�^�-���SE}}��mcz��褢+<�F�,��k�D�٣�%B��i��~v̈́�����������Dџ��#�P��M!�c��w3�<�6=��~�@!�q��L����p������H0�f��sY��@���������a�DSb'Xf���m8����'^����1X�ǩE=��R	�n�%��O�V��L��WDc���g!V��Ag��~��g s:�p�.#���}=������_��!�_��|E���ڨB`/o9�c�<�g��fD�.����O�p��ӿIZ�EF�]"��%�Fi�Lbc��"�Z��u��b��R��>@�����T}����E�(���n|��U� �
���GnW5�Y�,��A� #��G��|	���|�~�k�xG��T���� �j�VG��VB.�NW]*�Z�vF�s~.��T�<\�7�?��^z�|u��Tâ��(Oi�\�"�q�'�z�����
%����xe�I�wt���E�.^i�̾g�h�<�9�B4IN�;R��>�[�-���&h�$��U���'D2;I�,/<�_���vnkL���n���O���!M����H���S|�^�I�|�!~�q"YU�g�c��-{��(jݩ�R'�ͼ??TƲ�k9�~�hL$X�ڣLSRo5�u�����PB��Y���/V�"Ia ts��j㉜�{4��|qX%�z^U M��γ4�,��%C�s�j@5��~�� }u�8f�S��8�s0ǵ�F4��Ǖ�!�X���6=A��T�U[�X�l�.�eo���m��Ǌ�|@+����l	ݎ��xQBߠ!�S����T�m3l� ع;/P�]�'߽.�W �2��Et�`�L��݁4�ж�C�<�j��ڽ�x����HVG�w�HnȽ�:�ˎ&���_�/E'_�#]�����Ql�(ǚ��'���B�"7����T��V���hF�u��6�I��a,�aݎzT�By�c��e�=s�l$PTB�]��	���p�ׇ1ޤ<��C�ҭ�ܽ0c�����Q������j9��\/#�Ñ=�2��¦���X���@�'��(=}�[��:jiv�܁���۷��ψ_�/���*\ת~j	GW�< 0�8F���:ً�Xz�9m�$�4D��r�nx�ԫ Ř�=������׏q`��q� �A�]�h�\]��0��o4�#k��tQ��Rwdx���'&���Ѓ��3裺�ʂX�~Đ]z�.��Jd��!�-����d_��Ɂ��n�p���qt�C��g6)I���*i#fS8C��z1����wl!$(����@okDFE�r�9v�{~�,i@�ȗݤ���cv[*QT�0`�ր{j�p.��^��m"��P��@�0*S����D��:��n�|��Ǖ�c�V�������C��d���Xs�Ub3��Kk���{1�N!�N����'<��jΘ�r��9�v��c��8�֡����B�L���D
�l�>��[������	���"��+�7�ܴ�����%ׯ�?���*����\ZgLM>e��ƪA��L�c��Ǧ$�������ID���$�T�ǥMܕ�Q蔰G�_U�א�R�nz��kGy�T����2I>�1�N����;���c�IX�`N���C��.2�tGL���#�&c{_�]g��Oܻ0֠��~�{�s�A5Bh&x�SY@�Tt�,�a�FN����n��iz5~m��'�����q�h+��mHP<g����ԓO�.2!�&�͍˖|�@����yO��B�[te:�"�p��t �Zh�����ʺv ���C~��Swtx��
�L�9MI~��QW�T-���Ë�2���!ԡ?�� �G�|>P�*93OR�;�����=��- _���dy�'u��D�r��8�k��)��������@Zb����RZD���z�V�9U�� ���m�� SR_��7�����d�3E��p�U�b��y9[͛�?�(��s�d��̰E}wW!BQ��Λ�[�(�sC7�E���x�p� r��b�#�g�=̒��	��ᚕ���K[�}���_�J1�%�x2�V�4T΃i�X�m��/��j�&oՃd�?T�����e�C�v��BwHD���eCV�Q0h���q�ٯ~hi�F�}�r�؛��X�%����m���*#�I�Qu)�i�uN�\�9���y#~"$ׁJ1��w�KY�ᄅM�����
qmɈAYDF�	g�q�^��!i�
�Ar:��)@e^�˳*��{�
�@x��lw�	���%�W��\]9�?B]�[cV�tbc�H� �����d`�T�4�^�;B��Vj�+� �Б��Hcp�<g�����j$�͌�^����x�������w�2�b2*���K澄�n�U�o�e9�1�6h����^��ϱ��7�w���-��;�����B�Дz1�� �)!Dծ$	+�����T����|<����
���IF�]��g|�/G��`�w�b�#){�@#��$�u,�I��?B�_�N72�ԧ1��tN�|�x�&�� ֆs� T�T��:�%�k�l�
�����,V���������=o��4C���~�����4N��8�:ʞd���?t7��^�����l�n_򙛿��� EWx�6�P��<Ew��D ��$�"i{7����DF����������S�
�����x����z�.�0{J������]�e2ݽ3,z/��k4��E#����ݧ ��2A����;�lo�<�c����2/㈽*l7�uf37�Bg�T����e��_T�H��
��;Iu"@W��cP�5ۡ�b',o;���O��ܤ��'GQ���.K �,��o����B��Y��7}��!HG�fFL�"�+�kq"�.&B�_����͋C�d���u%bk�!/�5�#�"��QГ��N2�E&ѿ�2�h�^2O�ce���Qr\���~͉��	�g㾬�:�2ͨ1I5�n�hW��,o8 �O����eȊ���mۮ;xn���,��;00g��D"��=�Z?ޠ��O���q�����F���]��xS4崳|��M�b�m=�B/��Dp�)���O
��/u��<B�k0�5�4xO�g)��yqœ������#~9�,Z�0Lko�����9S��Q撾%|�z�;��j؍/z��A��`�v�m��P��P*mL�� �a���y~�~#��8z�	B��*_7�Y�¹4�!i9k�sa����#B�6ٗN!R�r�Y���}I]*O���C��@`��c�0SC�N�	Jm��,�8��"�U�ĩ'��qo�^���t��RɏZ�#p�8K��c�7�J���/�}��=��aOV;3�� ����6P"�z�烫���c�؈�P��B�Хq+�O;�����:S��lGW��XQ������[ g[�P���W�?��^1��s���E�Vb��u���'��?Z*i�{�"�\�:�BWs>��2q��� 5��V�Q0���'?�ݯH�����]��2���O�$>'����h�(�FQz|;Hɳ,�;�}~dfA��l��g��?����Bvs���e���$���4H��L�Y�CÈ4E�ʆ���v��Jդv��6�<ۆ	����Pau��~y�6)H�Z��|��d�T����e
��A���W
~g���Ѓ�H��pv}�񹈓gqo�t��E^�i2�k��Sd�I{S�-�S^YYR��b>�]��nl�%�$a�w�x���1.Y
Fv�����:��^������Y��xw�@?"�(�_�ݏu�)-q����id/���wt��츦���W�0�����ө���D�T�1��l��`\C�*1��[jѶ�J��;�:Y��a��O ҁ_�'���_3�W�煎�kl@u��%�7ҺT��W�w�L�����6�/�ɏO�4/�z��H���7�����F��ί�-ͽ!�V���G�e�Q�ҼO��J��\�x�):���������g;Q�r�mg
��f罆w~��5t> 0���Z�C;��尽3o�d���H �k�Etk5����
���y�7���{o���s뼕T���Du��g���˃��l\h�X�.� %�:����@�����^���x��xDK)[pn���8�|�GF�	�Ь���<��k�p�����Pɍm���uBL��.�~$c	���Y�	������$�F˩ ��sn�c��R�N(z <�LtV���bG�m. 2�En����8��d�|%�D �p/�e+p�"Լ؈�_G;�e�V�6'�YR�#|�N���~޲we��H��D#����7QI��]���hv��xi_q�L�����FǤNگ����b�3.����E�&@8{��� �R>V�t\t�UIo����`�{�$敫`�i6Jʅ1�	�{��o�W:�)�'%�A�.	}����Sf�zsѓ(����c�1l=ؘ�:{ZZ���bk�"UXx5�f�MYؒt����R���a��h�o��{�I����_��h�����Z8���ߟ��,�d�:�� c��a��l_��8`Ҿ'��� �;��s���=�3��Dˋ���{��.�Z��tɔ��j��d]5�2zvʻ�`�U����P ��N�$�t�*��*\��O�/�e\�ϳ�ۖ}ȮP$�4.�-�}��_�;A�osc���C�ڀ,�Xҙ�rBզA��ĳl��[-�l�+�����OܑK/S�E�K������ݡx�Vqd����m�Zʜ�W������ �N�Qo��|'��r����`?�X+TQ�� .�:a�ԇ!�zm{�k���z�ƪ
��U���ؕ'u����'��<�����X���r��9?��=Hҏ�v����s�(jp��耳�
l@���H�]�!���|j�O��6)Ա�駮h���׋`��mhλ@����ׁ��h�v��v%̻sB~�u�a+-�R�)���S�d:�����U��<]�H������f�x�.*�AzQ������c�?U7��]�3�2�ĸE Gg8ѹ�;�& ��c��k��;����o,=�*�tK��0��p������]Q�`���nZ�ȉ���ӧu�f���'1�]ʄ��������ڟ #x�'Q�Fe,|I��ܷ?�wuR��8W�.	��;*�;iami��RF��7%����=�[,aT갗v�dN����7�4{p�2]���W��p��,��<���:?%G���: a�v)�˿��:��8t��;�S�}u��QQ�����N�����%[��08DשfR�Ѥ]	8�>��U��A�يU{g�������^�z��J������&�i��r�J�pŜ�e��p��"d�M�V�O���(7�gV�������Q3�O�P��ӵ�����I�k|[%�(U��׽[���w��e�����d�#���]���i�&m4����P>�:t,�������YQv�VW�4PŘ�Ę��A��;:��������i��d�1�w�ք�GT �ʮ�_%�:G ��v:���($��z�֎���}pf�\a�K�6�OqIE���݁����L)yPA�'D�f�ʖ��8�.�c���{Ez�<biYٹ����Ԁb(�+/Gq�U7�4��f,N�t��(����S��w3r����2z
B��Y������=7hс���Q?�����P�����+��6� 2�)�	�1��	y$��;q��Y�*�Į���/2^�I�඼ϔ�S�w�O�aD
.����F�(���^������Z�#*?c��`Y\^�W���a6󔣪6W�������������w�[�|��h֛Q\���� g0W9�	�.�-+*�t�{�I�߀r ��*D��T�*�]a�X�H�/��g<��;UtX�P���=��-{W��Xz����6��r�t:��B�����qb˱Ƃ&ü+8Ԏ�m���R#gk�NT�6^�'��KS58'N��>W�}���q�݌�Ov|�<Y��e)�L��'�^%ENd����(�}R��ew7C����Z��C�1
��=H�{�v�J o�,���C��/�)�K��,��,17�]}B{0>�+�`���B�,�6ٔ/�+�m�W'�u����cѳ�$��.&[�R��6�N �@۠��,o�w��W(>���-n��A�r~U�b���
GX<T����^t�D-:�w�H�F��L�VcmZ�/n��U.x�d.��0��AB�L�� ���8M�\pNo�9C�O��wZ��Z��.�~��#��FL�2���k&�n�Y�u���@�J�r.�Fs���v��g��}�� ׌�����is�H�c���3�
�z{�W���� .z唺fr�"�.��8�{a�&Qe�>¼wq��1cB���ҡ��j���!� �_�RT�/�W����+�e�𫽆L�ï��^΁ꮶ���;>�lt�Z�d#�>�?�ʢ -����Sd_m>��TBz~�A\yo/>�,(���B���q��҇T�w�L�m�?��ӓ�}H\�L�n�i��翄-.S� ����;���엻+��L@_t�
�/x��/�'|�<�PuQ@�	2񧏧�ň�����(����h�x�8� �um��nrk��~�Ң��Ђ�?,�;.���u|�l��e�BH�ͷ�M�*E)���C�g�4'��эp:����e�%��P��vc����B�졉豋�K��\9����k�8W#���6�G1�	���^�X��,ow83{f*f�x-jwrlU�B�i�w��"�bl�sl��}��8\�+��ړ��ZG�NO� ��c������b��}4�^�20x޿�1�O��6V�� �����(�`��R�2��7ܳ^��>�挓eɔ~K�T��&��R�mĀ���'��J�<�+�<�wc+���E�7���K�Cf��6��w�I�����NFeI]�zM��j�wO�����<yڔ
�MEr��$1�`��V���0˗݀�(n^�q}7�I�m�T�D��:�z��&R�uc��z�����B��y�I���f�����r��4T���R]��;̔����B.A���/�O�Lx=�1���p�W#�Q�N0+� DǢ��R@�h���f4���,+�jIiV��`.�
qäl��J�:E�Y����M�I%ʹ��%65xR�y���Q2��)����;5>05�d�RA��/�
Q��ū���8rJAǊ�g�TQ��A.�-df0 'x{� ����9�@=�[��ba{�"���M!	6����
��3e�Rb��*x�Y7D�{����}�c��H[f�.[Gr�ߖ����;�M�rLe^u���ѷr���@�u�pW��O�,�I-��M��@a̱��D�2yZ$9h����F��}�:��姐�,�tA��3ٴ;�"�V%�Z<2���=��o�߱ N�w=_0���-���>��^&�3Ҷ"����dD��
�C����I���>�"��.�}A��<��mv��=��<_j�D��}���3|s��w� ���Č\�E(f�9#)8ҿ����b2N���d__f�i^������+t��bh���OUۜc�p�τr�Y(���G	Q`�dS�Ϋ�7�h)i�ȺA���'��8/���1�� 	�+� ]E͉�	bWAd�G�/C&�$l|��N�Y���ؽ�5�$\��r�*,p	QcQ���n��;"�b���T����Y�p>����mmEMz�Q�[�� uDp.�S\f�ΡLK87�Z���w�)����C<0��jbf��m�#J���{���(������u!�S��%�w�����Z|~ł�/J��b7D����y�*��)�cc��	�Ǒ��ƕ��?�gݚ~#� �&����O�~��2���l�:�aP"|j���ۓ�K=��q��Qo)�+�f�/�e������%�b��F���3�؋&k�Ƭߋy�i��{~&����x D��t�+����ѥ
��x��ٴP)�C�ZQS�ee�=_���Tv"ʕs�[!�LU��"�X~t2��@&�X�����V��gj5s����|���8m��PD1�;b��<<���H��z���ol��T�Bm):龸4g�y�ଌ���W�Ҿd;��a�.a�'Ұ���������4��k��_{n�׿�s�Pr��0���!%8���3�</�4��pfuD�)�.��X�v�ߠ͊��T�W?�YdPl�aY�x��-��0�jI"�������u��X-)j�e0�%�u���^��d@�����{��TW� ����K��	PL��Υq�ON���X�����8I��ߋE'����"]P����5#�AѰ�x�2������7f���M?�X$�z(|����hӸ�1��(�a�O��d�3*�5�T��٤LKD+�m#E��#P.gL�\H�ҟ��	jA������V��:c�����]>�_�.����w��q�2B����O��}�.�SAf��Y5�6w{?�sd��Z�%,�����ɄMj������(s�sȏ�Υ;��uvh�_k<�]�7z��j�~O�y���ǵ;�U�R���˱c��|dv³R��#
̧׳��4E\�����j���k�Y�����Ӧfr�+9|uu?��UX�6��%�O���|���Q8��8m��v�6H�/�ЁhXNmߜ�����U���͔������@�nw?�T!岨�'�#�ݩ�u�s�gl2p�*�  N�K��P�R��x/���1o�XCU���]2p7�Kϊj��@�0G�,@(����<��l6��m�?) H�y���3�6��5?���"}s��ى�-S���7�����a����i ���:$�i�ޜ<R���pC�q.���v@C��R���ִ�����
�w�u�5��P�K�h3W[�&(�!������Ƌq��C��DiƜt�گ���^:;�./���xW`��_|��L2�\ ,p	�03?����A����Bqc�B���?4�������-qϤ�2���(jr���e�[���{�� ��$1�&��o_S��ج���w���hkӝ��@CZ_W2P&U�?��!���D�w�.����!3x��J"���Z�N\�έ��?{>W����J�G:>�v)��)`q\K����[1��
`�G-Mv�Xf[�`��y�y��;����V�!�����%��[(D�5_ݺ���Ù�Z����.�-�llU�l��G�*�,&x$@�o(�����Y0���j��q=���t(��U|���lS�{@
��U���%���VC�Պ�Ә����3K�3}����.i$��GU�<��BWLJ1q��
�/��+'d4��	�"{l�ѣb�	��<3ݼ$�ON�&�̢7��l�;��ش�C�Z���n���K�z*��ZO5��(؊-�T��q� ps�W�+BS�Α�b؞J�Tj�ث7E��DEμ��P��!�ԧ�
�;�C��$�R�Ų~c^��]U8�YjF"��7)%��@�J��� x�ؙb�L�&C��M�
�G�LFʲ5D�M�GV����~�ouS�9�����r�ؤ�d�N,n���"tz1�C����X�x#H�|0��fthv��,"R���턓��Q�G3�mm1�L\�9$�h�)���%3�ڟ=_X代U�7��v��}ω7зb�.���\��ב�TLృ?�`��>Hsb�c��f�������Y�U(�$X�&�%8ry��Ëe+��,���-a�,��2�F ~%Y���D_{0��+�-�jp�a���x?�L���I�����HUֲc54�����S��_���*���1*��*�H];�L��5m=j��s%N�_�H�?�
����k�)	�&����`��ȁ,:.�<+>�G�Z�c�g���J���+��^�c^�A��KуxT^����Ev�v�i�d}�G��&C��O��#�ûk��[փm��!�Hw�R�p��>���)�u�r���QkŪ��.�x>fb��������*_�rv�;9ݞ���f{nSaMو�9H��[m����"�2��X�_ V5L�3�y"��dP�<1Nۅ$�
[l�GZٴ�b��4�Z: ��Ԩ��6ޖ�U �����������%vx�=:�+ Φk�N��f�_H�5��U����{��v��P� �%�,lz��n̳������Ђ�M��z�����?z�9��z%XG��Q��9���ׅt#+�c�y���+Hq�N�O���_�V��������,T�
G�e���+I n�WL�Fጒ�'a���F�"����S,��]+z�(��8�G�G�l˟�/�,$�TlL�k	3\Z�-h���D�H��iz%ܮ�������%�<�,��H�<�̒��.�["�	��C� �����o�J�48j��ܗ�����L���E��Bv����=8� ӻ��3�7cA=�]����T,L�'Ag�eb��>��6h�� �Rqeg7~nZ�G�?���Й����r0��6�Ի9Zz#���d�E�^w�:;W��S^X�.�܄lmf�x����Z��9C�Q�#���S��K��,]������HB��r��$�o��$�j�������_H����\1�3'�
~��1Iӯ�Jn��:�c�2O�V)c��%6�7$I��6D�2�5#���r�)�u1Nvk�%7K3	+l!J�q/���ȼ|\R}x�	�T�k����ez��Q�&�P,�+��,��6�����)�ɴ���W�s�/(�CjuϹ��^ީ�֏�����Es�e�C_�����)s�gw	�⓫z*�&���#����1z�vM\�ǌ�p&����H�Rg	6m,9S{׾&�?����"�ʵ���$��3&�6�=$�v�o+ϥ��G�zI�C\2�Q�����`d����1�c/0��̧���*~Ǿu@ 9s�E��͖��w�d��c��2��&�AsD��r\Ґ+A� O���k��{'��_3E��`"�ssܸ��{ӡb�$�f/�S~��SX\_�����cd?/�/���葴Gm>�a��}i��<��l5��HIW *�C^�|���O�ڀ��ǻ!�6Eo�9j�cXeaM>�*d-����AyJiM�M�DG�l��w7r����n?��HT)����e۰Tg=���V#���\G���d�r��҆�YT�UK��V�|`�^A��W�Um���B0H�������ճ��pZpz�l!�	�9�n�ϔʥ�S�����Ϊ���M),�'��SKH�[�}�&Ct��&�$��0���_��i3���ؾ�i�z�T���:*���x����h{冸��	�}
�Ѝ�L����6�@j��*�P��g@{jI�Ȝλ���^��>�kb�7St���)��
�BT�Eeۆ���e2�����h	�QnZ�rRF�#3����`�1HB�mkrڹ̳�Y�<"��k��[}u�`gV|�V|Ջ�a��QQk�F���)�[��5/ݦ�R w����Nz����K� 3-��4��HUG�>߈��'�"X�x|I��� �i�;���I�W�t��u����&S���O�xą�A������(�9���J]��	\<a��=wgЦ[�Of��qiC�ȫLoEh~����˪O�Mھ�;�TTBvR1������s|~1�����\���/8"�8smU9�l����Z�C&���śupm�g#.c�b�D�R��l�g����B��>��DKbG�R��%M#��B�~[�:݅��b�׿�*�
L�xwQ�`*m̏�����Q�r��*�L���*�����Y��Nw�嗎Lґ���͈�KQ4uX�2a���ƮR�Ggh���A�6���|�E�*8�A�fY[��B��8�:�AX�;x���ӫ��7�(��	�-��F��>K���2���+4o-�c�H�R�L�:�%��~Z�ւ�}Q0	�#0�yv�n�1�MCX��iU��5gm%�<R{�mn2��-�0�s�9Hd=����y�t`W	H���I��N&8WBV xH���=��К=&I�;aF��հ]�
����i����]��5�i�g FB���c���(�{��QB��H�l8a��y��.-h�ET��2c�U>e��G��Q�b���{%:�eh>HN��s-�xz�3H�����'���.�ot�t�-9p�g��ad>��j�E�u�	�֏Z���G����]��@	bܽW���6SM�ݵ�Hݤ���0>���@I�&�����(%����]e�[�T�<���%���=���IArï�{Ve��S�Z��	F�C���'ӥb�
-�e�4��?I�U�š	�G�(�W�̆�>P�k�I��7U`g:��<0>(�Ƴ5�b����L��
iէ2ŏW��qUV���O#��v.��������i�Ԗ��.�P?�6��u�j+='�A�MV���R>[8"$'[����J�'hϙ��I����;��Ʈu�䭬��Py�}s�R?�*��&r��r8*)��@H����(gp�#�6�o���]�x⩣Y	�Q�����x�R/B�������y\0�>fr����m����L+a��_�plV�vhF�ҡ�S`���Y\QKdt8�C3�GT�:ž4�Q�Zd������m��n�z��q�\+��.���G`-���仺,�>W:^��_W�a�QUC�3-r�5W�Kl�
��zV�M'�v*�k=�Q
�h2���+)�#�B�o���&���מM�b �3�qOzed��\����^��~�yR��\�|u��^�:��c�h��Z���֩�H��y��Bm���{\#�wY�ڣ��Uh�%�X��ӂ��dL�Ag����ov�����w^+��p�5�m�qz�l!���w�P@o�(����?@��-�!Q_��/~��C-Ml��Nc�L�0ض�U�ϥ�����r��E��}�I�����%πDm���Q2�?�$iwqɻ�H��2��vz������3v�����$o����p6�W^�^��nOi�}��6��m��5����?)���~��̖�}���#,�w>ǩ^��O��da���D:��cjq��V�}�r�k�7T�qa�Q{�/j��[��)].�8n�*A�r�Uu�����޿k��X��}�fed�S�h�U�yu��*�!~��ªf@�e!i�pu�R��n ���0�_(\��>W�E�J>�7=oF����bj$2�a���h�h8��	�\�h�<�"T��@�<�OD���>;�/"Э(���C�7�QL|hh���8AY�e��^ë�|�+����Z1��t˅!�q�&޾����L�
��4��Z�rR�@3Ν0�z������7�B��G)�%N����I$Z�Ʃ�-��Λ���NL��f���U�Ȝ|k*ot�t"���<�E�\��hǩa� ��;Sl��4�'Կ-�\���W6 �z������m�-����w��\hP 4-4��
���xf���A��}8UO|C����%��4��I�b��TهjXx���*��@����`%s����H%��n���?��oc<��?޵IIl��6�{H '�Ba?Qu	�jH���16Uv�s�1��O%���u���q�1���w�<�v%fY�~�&���GiǦ�I����� 4�[u�#7������Ic�S,��^)b��}z>g� ���x�����'�����HH,�ւ�e��5�.�@��$Y��q%v�Q��RW�*"4M�ʂ�s�#Й�iתm�h�0^{���gPb{$XN�)}og����&��0zy�l/�ψY�S>���A�[E|¿{��rk�
�ה�(O���u+�O7�Xc����.l�҅��
jsA�<}\��2j����
�����5M��F�Ι��ٔ1�򻭢��|������3���,>O�P�٫e�P��#N86�,(�E�lS�G�ͯf��Y�|]��ɾ�.T��/4�9Ķ�&N�|=
��B� �el�� �y��M��f�̀����@Y�	Oީ�X ���sWA����P�ٍX&K�"e���l:K��^h�PE&[8��쑭҃x4���l�NMH0y������ �� ���>�6��Py���Ґ��#����{GD<����ٰu�'�"l��4g��	|y|�w���9�l����:�9s׌�iص�L�MO"��/GW������^�wރ~�&���}�7���"��)�z+Ca��lvO��+).�q�b�Y ���B�z���_�\s ���v�j�]�-���5C�r�@I�y-/�kI���ۗL�
Jq?6Ҏ?��ŋ��8W��*8���=�}0y9��q�m�3��l^�a���՗`�S։䪑��';E�#�I��6�}o���l�$��p����J
3n��Oe��̓��R��S���΋��ӹ��8{C�yLƮ���f+�:��&�7��lK����SqMH4@� 0�Ley�p(�*��]~�� 4��.FϬ��������������)�Ϟ�$�T�N���������TK�9�U�5����]	���β���O�H4�G/R�>��+�(�ɒ�)�S~P��t.na-F+V|P�	�ms�l`XK8��O�ƍ�z:4Ή�ʜ�8�o�2��B�1�ڷ=�w�lKR#�&��ӶF��b��WX�Ğ��er6}r���������𷄲��Z�)�[��ٌ��R6�����2i,w���\�p����]���bB;��������J��\�s��KNz���d�*��!ۄ$Vuvqc#\SAv*�\)胇k:����[� ]x�����6�Y�byj�o�݈]���҈��v���%�<.�_Y��+(��JӾc���[��K��������ټ�_`��^�;B �VڠD�ϖ�ʴm]>�s삳&��r�mT�?J+�ml�?b_���
�B��
���L�9tS	Fm��hiAVtk��2��J� #���g�t�p|eI6<ww�x��ɍ�`$�P�'誱�V٥�H����x0?��5׶�ⴴ*Y�@�y��񭇷d�����!��v��X���;n_����E���f>��l񝶿��j9Uj��t�X�{������kȻ,4+l�%�h��t���6g�!��Ƌ9
�S��a���Lc_��I.f��(��$�,��c�y��fA�t��v����~G=<s�~���z��{TH�IԪ�ȭd�P3�</F�e��u��k�U�pL���g�#��$�+Vx�3��hy����
3�'�+���$(�6�V�3E�0�ɤ�]Cv1�Ѓ{z5���1�z��ېⱧ��d~6���ƇN�L6׈��a㙌>Q ��r�@k������*��ÿ]��8(Ẵ?�4+a�2�pN"K2ޤ#ڤ�\3?��;���\c��g�	�B���1h���t�&Ȫ���2���Q��x���(���-�ZWB��T�ݺ�����̺�K����ʤ����y�=�q�����]"9&����&�˭ʤ����ڪ�����,�C$�b�� ��j��¥A� �C|�m�q�	�T^�}W�ʵ_Ɩ�0�3�����aO�������{��a��i��H�5(���i�>���4���|Y��u����Ys`<I�^�Ķ����=l�`�ڂ'p��Y�D�9H0���n��33fD��<_�,�d�0�_���/�#=���n~�%���K�}�@��|`�C��X��d�Įc'(���qos��=�n��`Ok`[wE���6�9@o�|]!��14H�O̪�t�� ��*�p����}�	��-�	A�����VT���ܑgV~���<�EA�������)Hg]�&����K�8B��#�B<�����nI���A��n�1���Z`��as�I���R�:��[U���W�r�y��/�z�\�?�K�ёQ�>��F�}������z����wD�pތwTO)*��S��'�5�����,����(@���tdd�ȓW��|k�d��֗&{�fQ�F�)�nܑ�4�H%MAA���
��n�'3=X�}YR�XB�6nU�U:T����:�3�����EE���'�x>�;�!f�JnLv��K�;��_\��u��m��Z�-�C�O�F�$^��Z��qX�&���Q{)�<���<�|�C���{dIO�p僪/mmS�ٿ�F���b�>��o�W�?:ɵ�m�A2���0�dT1G[���)fV;��FP+{K���J�_�OG/z�� 4]�<�����CT��0|,:i�dm�`�q�G���瞩P�o:��z��-³jJa��=�f�g��
�:tѭJ��q�ڦ�)<n�4�ȱ�v1������;��7���������N�wk�ߦ-�c��<L�4O5�}*h�Ci,($���y��3���WN�g�࣎g�"ڛ:P0�=�U�Z���D3l	D$�9$��XW�`uJ%�P5� ��������CA��a#i� *��s>6��`�)+��W�K5wX��� �ny
F����h��/p����X���b���}bm���V\	��r�=n�.����)c�}KpO�$���$�ݞ&�e�T��y&��o�Rm�������4�=����Mcs�I�g��_|&F��������$�.m�Ȇl���C��k��Xh���3�xL6J�/��/?���y6 c�iC�������1#����"[T�l�P�!H ���dV�@�d�
���[���Ջ�'q'"���x&� R��`�Q�6�'�� ��R�f�K��{���sEI��hx���]�o���2M�Q>Ĭ�cY.��6$��$0Ѧ��^���K�G��q��W]�!��;=a�E��N��[��.�ˈ�*Y��Z���"g�b1gWUL��ؽml�y�Ut4N�׻�n0��-O�����.�c�\�����.u0����רi�3J�;��Y���#�B���a��;����1��}H��	M��Z�>#�lc>V�EHS8&`p�R��:2>�}�ç��i���,��u?�L�S���,Dwi�n��ks	��N�ξ�����7$�̈���MC��<��Q0�t��(Pl��C�8�Ah�������;P!Eu��,�N�R_)Z#o��ˇ�=xi�o��R���>|�Zz4����2��G��sv�B�F�m���Ƣ\�+��<@I0��p���>��ޞ�[�"\�8ŅϠв�����L%��F��
�p&a��]���
��ɷ�w�y^d`���_/+S�V}�(������9WV�մVh𲅿<}�9�P��Ru��m^�~k�zl旹�]��Ƶg�fG��9�.>���O��e��$�1�8#4^���ԾH�iAw�A���y�����Ś�жP�%/`�	����*�%�+k���=�7������Txw!)�*�Z+6�#:� ��@2"�T������o�o��i Rh�\ށ�i�*�<;���0LH� 4�"?��I=�v13qs�Op��l                                                                                                   