MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                       PE  L 7R�H        �            1      P    @                      �                                        �  d    �  �                                                                                                          .text   �0                          `.data   �Q   P   N                 @  @.rsrc       �      h              @  @.idata  �   �      n              @  �                                                                                                                                                                                                                                                                                                                                                                                                                        �d$2�d$Ѝd$�v$��  ���D$��  �      $�  �d$t�d$��d$��$$  �i
  �d$-�d$Սd$f� ��  �d$r�d$��d$��32 �;  �d$�d$�d$0�8  �d$	�d$��d$hF\��$1$3�$�d$[�d$��d$�  �d$z�d$��d$�d$��$�  �d$�d$��d$�D$�  �d$.�d$ԍd$�t$@�  �d$f�d$��d$�d$��$�4$��  �d$z�d$��d$�<$�d$F�d$��d$��  �d$?�d$Íd$����  �d$(�d$ڍd$h��C�$�"ʑ�$�  �d$Z�d$��d$hq�fz�$1$3�$�d$F�d$��d$�  �d$@�d$d$���� 
  �d$W�d$��d$�T�  �d$y�d$��d$P�4$3���p������xIg�4$�)  �d$%�d$ݍd$�d$��$�   �d$�d$��d$�t$8�3
  �d$�d$��d$h���*�4$�GG��$�  �d$_�d$��d$f5��h  �d$b�d$��d$v<�  �d$u�d$��d$�� P  ��  �d$.�d$ԍd$�T$�	  �d$E�d$��d$h�>&I�4$$3�4$�d$8�d$ʍd$�G����d$A�d$��d$�d$��4$$�4$�d$v�d$��d$�����d$�d$�d$����  ���d$O�d$��  �    $�    �  �d$1�d$эd$ho,�j�$GU���$��  �d$�d$��d$�@4��  �d$�d$��d$�L4�}  �d$r�d$��d$h��9�$1$3�$�d$t�d$��d$�,  �d$H�d$��d$��{-��{��
  �d$Z�d$��d$+���  �d$0�d$ҍd$W�$1$3�$�d$�d$��d$�  �d$�d$�d$���7  �d$D�d$��d$���  ���D$��B����       ����d$\�d$��d$�d$�V��h�6'`�F^�,$L����  �d$0�d$ҍd$�@�����d$+�d$׍d$�6�  �d$d�d$��d$���F   ���D$��  �    � &  �d$^�d$��d$T��  �d$�d$�d$V14$^�    �����d$`�d$��d$V14$^V$^�y  �d$�d$��d$�v��  �d$\�d$��d$V14$^�   �%  �d$y�d$��d$��"  �E  �d$+�d$׍d$f3��  �d$"�d$��d$��|�  �d$v�d$��d$��$   ��  �d$B�d$��d$�d$��d$��$��h�<N6�4$�]"f�C�$�d$I�d$��d$�  �d$�d$�d$�d$��$�$�$$�����$3�$�d$�d$�d$�5����d$y�d$��d$H��  �d$�d$��d$���j����d$5�d$͍d$f�V�&  �d$n�d$��d$���  �d$#�d$ߍd$W1<$_W4$_������d$8�d$ʍd$h�f!-�$�~L,hAE;1�,$��R��^j�$�E�,$�d$\�d$��d$�  �d$u�d$��d$�D������d$�d$��d$��  �   ���d$-�d$��1
  �����d$'�d$ۍd$��   �=  ���D$��>  �#����d$R�d$��d$��$�����d$S�d$��d$QS��h���'�C[�<$��   �d$f�d$��d$��  �d$t�d$��d$hI��)�$�$@   �����d$/�d$Ӎd$���=����d$g�d$��d$��$  ������d$#�d$ߍd$f3������d$6�d$̍d$��    �	�'  �d$�d$�d$�T4�  �d$w�d$��d$�$�d$w�d$��d$�'  �d$�d$�d$�v`�b  �d$W�d$��d$�4�+�+�+�+���  �d$N�d$��d$S1$[S$[�����d$9�d$ɍd$�$��  �d$W�d$��d$�@�	  �d$x�d$��d$;��   ���d$1�d$��  ��	  ���d$�d$��*���������d$�d$��d$���  �d$K�d$��d$VhU�cVh�U��D$�Т�d$�,$�  �d$F�d$��d$1L$(�����d$z�d$��d$d�@/�~	  �d$I�d$��d$WS��h���>�C[�<$�  ���D$����������d$#�d$ߍd$����*
  �d$v�d$��d$���]  �V������D$��;  �����d$I�d$��d$V14$^4$�d$b�d$��d$�V����d$�d$�d$���   �d$�d$ �d$�$�d$5�d$͍d$�%����d$+�d$׍d$U�$1$3�$�d$s�d$��d$�����d$#�d$ߍd$U�$4$�$�d$C�d$��d$��  ���d$F�d$���  �����d$R�d$��d$�L$�����d$8�d$ʍd$V14$^V1$^�  �d$n�d$��d$R�4$14$3�4$�d$b�d$��d$�  ���D$�����������d$%�d$ݍd$��$(  �  �d$G�d$��d$R�4$14$3�4$�d$K�d$��d$�����d$B�d$��d$-   �|  �d$�d$�d$Q�$�@绉4$������d$�d$�d$�L4�����d$O�d$��d$Q�$4$�4$�d$�d$�d$�  ���d$I�d$�������  �d$V�d$��d$�d$��$1$�$�d$8�d$ʍd$�����d$�d$��d$R�$�$�ꔷ�  �d$!�d$�d$=   ������d$ �d$�d$�4$�d$�d$�d$�K����d$/�d$Ӎd$U�4$$�$�d$x�d$��d$�����d$�d$�d$��1  �d$(�d$ڍd$W�$$3�$�d$I�d$��d$�V����d$6�d$̍d$�������d$�d$��d$P�,$1,$3�,$�d$�d$�d$�D   �d$g�d$��d$Q�4$$3�$�d$O�d$��d$��   �d$f�d$��d$P1$XP14$X�����d$L�d$��d$�d$�P��h���@X�$�  �d$B�d$��d$�v �����d$:�d$ȍd$���>����d$�d$��d$���@����d$O�d$��d$�L��  �d$�d$��d$S�4$$�4$�d$@�d$d$�����d$�d$�d$�6�������D$������    �  U����d$�d$�d$R�$$�$�d$6�d$̍d$�?����d$�d$��d$h?�}	Q��h/HޏAYh��,�,$��RP��h�M  �@X�E�,$�d$a�d$��d$�  �d$c�d$��d$B�M����d$�d$�d$h��J�$g!e&U�$��W�$rote�C3�$�d$k�d$��d$�����d$6�d$̍d$��� ����d$�d$��d$�d$��<$�$Virt�����d$O�d$��d$�T4�����d$[�d$��d$����   �d$i�d$��d$T�������D$��?����P����d$O�d$��d$E�2����d$T�d$��d$��$$  �l����d$>�d$čd$��a  �d$X�d$��d$�T������d$�d$�d$�2�7-�2�7�(  �d$��$1$�$�d$M�d$��d$�����d$N�d$��d$�L�
����d$k�d$��d$�L�   ���d$�d$�����������d$g�d$��d$�d$��,$�����d$#�d$ߍd$M�����d$L�d$��d$A�����d$[�d$��d$�T,������d$p�d$��d$�L,�r����d$3�d$ύd$�T4�t   �d$w�d$��d$��������d$;�d$Ǎd$�$�d$P�d$��d$�,����d$�d$�d$�����AA���   �d$3�d$ύd$�������d$(�d$ڍd$������d$p�d$��d$�T�����d$g�d$��d$d�@0�  �d$/�d$Ӎd$W1<$_<$�d$U�d$��d$�Q����d$^�d$��d$M�����d$,�d$֍d$S�$1$3�$�d$
�d$��d$�����d$=�d$ōd$�d$��$1$3�$�d$r�d$��d$�����d$�d$ �d$+W��  �d$@�d$d$T�L����d$�d$�d$�|$�����d$�d$�d$3��   ������d$w�d$��d$RS��h��掏C[�$������d$�d$��d$h�;Iu�,$�;Iu3�$�d$	�d$��d$�7����d$*�d$؍d$�������d$=�d$ōd$�|$�����d$4�d$΍d$��  �����d$&�d$܍d$�������d$�d$�d$�������d$�d$�d$VR��hu\��BZ�$�"I�����d$C�d$��d$�L4�����d$X�d$��d$�������d$�d$�d$V14$^	������d$i�d$��d$f=�J�9   �d$.�d$ԍd$G������d$d�d$��d$R�$$�$�d$=�d$ōd$�������D$������������d$\�d$��d$U1,$],$�d$I�d$��d$������d$�d$�d$B�����d$e�d$��d$h��W�$�4$������d$M�d$��d$�@<������d$D�d$��d$Q�$�$�$$   <�$3�$�d$<�d$ƍd$������d$(�d$ڍd$UWVQh�2�/Ph4Eh}�:2hS*) h�9��D$$��ލd$$�$�!������d$k�d$��d$h~Bщ$�$������d$7�d$ˍd$�d$��4$$�4$�d$1�d$эd$������d$$�d$ލd$V14$^4$�d$Q�d$��d$����                                                                                                                                                                                                                                                                                                                                                                                                                                                  1�Z�n�+��C���L'�}d�W����r����t��9c���	�ş���W"�OSo���=�C����K�����X�����{C7T���V�I�����$��W�������	JS����,f�$~fu2�KX�nAͼ��Z�4�$��}���k������L�E���x�x@\T#+<Sf��O�N$z}����u��D
/mm�7��t�>k�:��@��K@|_�'��I�{����L��f�q��Z�
�)��D�9�_�e9��*0-��e캪�cտ���8��HفD���C'[Js�	��,ş��'c���}E��:N����Z��J�YP����c��%��֩!�A�.�T�/j��0����\������;�V�~�~��,I�zj����ʚ��Ћ��o��ޜ*bo%��o�1x/V��K-�x�j�`V�o{�e��v�m�1�e��{����e�´c*�<7)��ي�B��J�U�� z����qї��E��A!�kr(���*�(;õ92�L����$,Μ�v�P����FN~�+�KZ\�Ԏ�7(�c�JW��ߡT̵�#��/�x'/p<�7�5*���̏��I�u�j�����4�[���z�E�������s���Q.R`;����a\��'�@���QԲ�������2�0�r��9e�����}(-����O��8��F�4k�h��Y�v�I
���BɖŰ� �)-�S~ܝg=�������	�w��P�g�G�'݋BIN��l��xP�>�,_̀��	�h�bØ��������5%���1?3;D����	�6��Y�һ8@R���S0&Z҃���$�������<���Ći=q��g\4J�;s�� �+�:{i���G�E��� �J���D��E�p��d��H�T�Mi��H�$�k��M�B�J/�6�vʰ�~<���G�����Ä���^��������A�JfQEmg7���"�>j����}�౾]4����9N�� �����3���㫌v�2M��QQ*" M���"��ٮ@�E=���[�֏@�8 �ƪ�'e�X	�+�Nj�ԗ�]p��?�oj���<��]jƌM9�M��;���O��7+m�]^l�4��� -��1,���߳��ALD�,R��&d���C�JTsCQ�Sɨw���nj�ԩ4u�<*������`�ȇ����b�a%��S��NX*�B Qd�X%��
9 "D�,͡<��U��L��m/���E_�:��� z]��k��[u}��aO�ac'�,($3�$*Q0N���i/$ekuw4���Gk�b;�7HZ�t�w�S�S� A�DdIe_����d�,	�mTФn�HW5�TQ���f����E��<ƥ��f�քB�{ۈ�chs%�g}��Tn��TPE�L���M�W6"L�)R_8��/�]�"-���Ld�nt� |%�XyJd�1ޝ�M�{Qi[D9�f1�פ��c�"œF��;����]�4�v4"�J|E	U�x�� uMgf��H��v�w���{��S��y��~p�
N�񃎦�,��l�M}<9 Z��{hض���V͊���̈́�u�Ĥ� �5n���P���A��}�($�-���=�O9\��`)V�Lh2b6^�Yxv�u�����HOiaؒ�5��Ho��`qrM�*:��#rTP�����i�gl:��Vm�m��´��¿��<x2.%�@
�;�\I�d)>p�}�/K��@�.|
�3^F*0F���:����3�0T�V��(�x~ܣ;�Q^��u��~J��>�U�UԔ"2�k-{�|�71DE����}ȁ�%�����}"�u���ّyJ�F�}�����{_��NИ���+=��|8C��\�O�_��9m��F~���uwazs�IS�r,'N�&�`o~�Y:F���w�1��Ŗ8B��^2	�p��v�����u��Q�⛦�2l��P��ҥ�V�_-	���!�3F��Վ^+d}����t�2�2^~���H���Q1�#6׻
��<�{�
�K�1�oާŁ5�x��@5y�M��#��os�h]�̂-�������R�幡k���y�袈�ƪ0�񟀿ÙC��[�^T��-��������&@���&5S7Z^��?8��ݰ�*���̝���Pֵy�:2���Fjj���A��f������,�"��q�#�^ER����U�ީS�'r���_�h�dRuX4��I�Cw��0~U=��P�`qR�
�KE񑓵��7����*"��k3د#��V�|=��es$��EH�6v<���E��6JbG����~g�6����U��^��p��*K�f;�fY��y6.������A>�F�6� T��0�O��{q�)���>7u/+&�4��C�e�9�쉷Rķ��u]�U�����Oܶ� �����?��O���"��L����z�:��#��-Φ$RW��|>�e��hʏy�+e��r�(gb�i9B�BwtW�	o��WI�J�P6^DVȘ'1��\�~h�y��H���;���){^�&uQa8~O��S�6b}�$r��Ⱥ�st��w�R��G$D3AI�$�V��cl|e�>l/�6�t�S����� �`��E\�����P���VI���*�]���\ϹndcE-�.�[`�n͋���P!�Y�6^/7谅��5-�UF~�G�t���������v��W�����W�>*�q��3T$* �WH��>4}㐷����3+����J65m��0�����q�V8@ө���;T�>c�⚆UT�>� �.J����o���\`�,@���ky���PL ���<�,T���G�|Q����|,R�ƭ4����њ\�KT�K
O)C�����E� �=h|���O�I!�Yp�<k@� r9��t��=@���Ǹ"���N�yD�SX��j�(�a�њ���Լl�Q9,��B�xeV�>e��a�x%:
��1�xJn�_)�'�~'�>Tx�ޘ�1+�95�T�x�ׂ�jN���8��-^r2z�[��G�_�)�1i�ڨo	Q����&H��)����V �z� f�]��OF��ATr}aՂr�\� ��*�-���N������F��M���PP���ԤO���:�jW��F*ٵf�,�_�s�[�6;�)����4�(��e*z�A�@-�}k{��E��dl-�c�%("c_�2�N�6� �md-&<_X�2yϜQ�U	h�l��x��k;b�-�~�/���vۂ�})��N��a���`�"?����q�ɭ4�)�[�W�=f��F�v�׬�gU A�e.1����K�h��b��}�j��
��γ�����/�Ѻ `��*>��� h�e��tz�>0�}�)+�!�\�i��KG��1;�)�vty*5Դ0o����Lk331��D�¼:^9�,'��F<8~�FTJI���k��K���5�8K9r�wq�"9Y�jbL�M��~d���BV%D%��T��_��
.�ԃsl�?���%G1�~�߻�=�^��􄋇�L��Բ*
��{z��=�V�����a��T�rn����p�Q�d@��S��ț`a��{���[�OW�䰸y�2�&�E�#��K��rug}l��C0u��Ep�m�6O�e}��"=����EZ�Zz�b+;�N��)S�cK<{*�X����e 78�v}���d�	Q��M\9p`�I�H�S!�����$�l��v�����J��~���=g�
캜7�~;j]i�7�TM�H���Qa����x��Y�'(��X���bhWp�9��%�=������ 5t���:͋[]��̮L0*2�ګ�2J*[<�`fZ�P2o��S՞�a����+��{{'���5q}VP�s�Y�}h�e9Ww;"�\�����s-�C���W���K��7�y`N����7<���Kz2K�%]�*��k���S�iw�dXE�-�&��v2J�u��A��eb�U�`Tݯy�j}��y�춅����;s����{�hW@�z�9��b���Ġ�~mDe}�L�ʁ���wm��t��������engؕ{�W��-�V���C�	e�����RtMx7<��
��Dl�C��$٬Q]�����l�oTP �R1�Af'ٳ �Z����Ԓ�+�F|�cq����@���,E`=�/8+�o�߮��c15�]�zPRQ{4H���D�
 �e�u.��B�lP�tN�%�n�3C�^�1c%i����<�F�pG��R�HB`��]n�i�Y��D���۞�3��d�aN+f}�-%9KG������bҁzC�>Y���߃%���Y2RiuY
r2��u
��F���rj�\��/�єiE�I9s�v��,��xJ�hf��{o���2ݠ!F=��wׅ��f�,�J9�%]�Cn�����+�]mZǗ���咽]LDN�������!�� &�i��2��%��8���� �=��J���׶C�S�G�r)�LQ�[PE>o�t!�2M�ߛIWd��Л^����;-�> 2�!,�""��^i|j��ئ��2�̃��+�:�G�T�枬��H�#F
������r8��d�Nl��cC��(�����(L_�����6�U"3<�+n��	|�E��_�)p>،Ug�}��"x�ʢl�q~�h�6�h�RV7,��[�F�� 8�O8�^� ߈�f`+ʈ��9������:To��]��#�5i�ͦ�������G��~t�X����!!��qYcB��t̘PNd$n����r8ހ���q��{�H��� e�>��lst�PGfwF�^ݣj�
B׳@�����[1t�.aZ�n?����-���`���Έ"ᑝ����ƘU4��m�\��\��wܨs�"���Ŵ3,\�[Ŋ�й'���Q2rz�O��������}�q����.]���;�&xZu�5�_���W��%}1aΙM��$�	 I��f�R� ��wok�H�p.�}J;p4]�ej�u%�Py�o�Qϙ��'>��8:Hr����/-z��:�Z�X��1���Kk`�zא� ���2Ix���f{l���d���I��d�d^c]�z�b��}��I'����Ly�eK��U���VjP�MvU��iUPV,u��V�Z�L���ӘZ�[ ��1��쾻�
����������H�/SR:��ֹ;͈;v�N�kÝE���,�_�S�I^4�X`�-�e�1���:�֝b�t��&�o�n� ,%s�#V����#,1��?(�i����^[W�y"�E�	���7pp!f��%Fl���w��v~b�Gc��L�~�_-D�B'Z��ڧ����[��dF$��0����	lm���	���6�Լ�R*�ң���i�U���S $��5�s��R3%� {����]+�*_�Ѕ�^�����EWȡ��n8���*ڥI�N :6�q�aAT�#c6;��k��C��L�����a^��?�����g�*��w���3�I%��E�#��ת��t�|_���*����dt��!"�<PW�I���"�evSmG��^�Ɨ�7���p̒�A�u�zd��+\L��ZZ�� ���X�=� ��`c�z��� �~d�C6���-{c�D�(��R�e��+*�ErI�h���z�l�*pM$��%�G�hD��,n���F�O
9튖$�
f���7�eO$���j���d��wMuO�y� 4�_\�a7��RԴ�]H������l��)ԟ�N-c��v2�_?��50tv�*�5����I�%�ݣ-���6�~��D�y��lJ����t<2h)�,�Wi���*��l��@�"QsB��[�����]Ƽ�.�>�/�@s[t�aǸȗ��0՚���+D��J��Yg�6E���� ���G�"gѲ��}^߾ڒ����۔Зd�:vb����Zj}�o�D	�f�$gE�+ի���R00��}�F����M�g3���,lm��뱀��|rC�V�Uw�U�d9���r9;�Uc��������}�`)��M@�O�������1+��F�K��7Śm�����2U�ࢯܾ��u�
|���E�i��:k���;7��Ӑ�w���b�����.�]�њ�!r�����-�g����T��KE��A��=��he�Ef�{����K=�B;�?�0��`ddAZ��y�C;T���@��R[�;]	�14����H��}?q�9�U`��uP�7�LƔ�g�4m)�dY�G�U�U(7N+�9��E��/W�DF	���[�*�N��*$��3&�oA�L�`��{)�ޡ߸������>��;@;W�_�~S;���(��
:��M�BYU�����x���N$�J��t���7���s���x�o�^����З�a��F�b�8Z�t;���2��25�'{+�L������ҢRr�H/Z����1~��2y�!����"��I)`��T�v�x�n�$:���9�V�!�z����$��gWT{G%k%k��U��r���4G��Kޞ0N}��F&��.��"��$>ԛw�_H���|�qP��S�W����	�%��$��nYw̫��7g���IDk�·-������a�"�bf�*�%%Z���R��Ȭ����#��׮A�B/�<�,���,K��� ��}
s@�8���7��a�飄e^D�[+g�ti��z�B0��p%PH�����:��a�Ah�t���n�;O�wW�w�����JĜ_5"lD8�k7Z�3��Y�,�M`�����&5���M���PnǕÌj�i����F�AT`+��[���At?Z�W7�^�j�$�Sh|����[cn��o���"�͊Pp/�u�? C7�ް���-�%e�Ǭ!��@H���tѳ�����oe��ˣ�H��*�C���@ٕc�rb�z��Ɲ�Mz�ݮ�����|�y��p��Lcw��PѥypU��R��z;��:b�}-
�͘�w[�tP���|���M)�b�Jĭ����P���w<�^�-���]ę��oC�Na�7���[��;ᕷ�q^$Cp���{��˶�Iy���;#^Wd�5�晎
��M3��ѓ��;NҧQ��;FR`w�t_�F�^�_��ꃋg�uf��w�o��B"u�f�	��
Ɨ�b�bD�kf�
�����k4:e�޲��p����f�:B��&<@�u��׺O��?�pmľsv��d��Q�+�}T�ry/�F/Ak�F�[P׫h�C��I��U}����
v�l��d���N�L�\\��㴃���f��zX����/]r=�xW�$KOu=ֲ����4��s�lUn��H^᳡��'ǟt��LF&[>���T�Ȱo���4k�@�anm�[��Sr���Y������n���Y(U��Bх���#F��VD�	-�%ӗ�<�� ��8�a�i�y�95�zL:�:+��-���ȐO�e(��GEp��g���RN�� ����B�G��H����5P�9珝�T&�*��J�~|�g	0�D ��4RG����U\i���t���	� �<�5�6$ ��NV��b��Fd1����;[a�=�O�a}M��f��xw\�8�	T7��ƴ��G4P��! }����Ӄy�L���1d�#౽�@�	I�wQ��;���(^}����J�A�9��(�?�
O�o"X8�Zi��L-�w��A$ �^�l�"�����	4��ޮ�B�4�K�jF,eEW�m9פwk��K�]�����o��������{w�*e՚F۩!�f�L)f	��TI���Ⱥ9X+Fg3�),!:>�6�х�NV��Z%Ls�x�0��Kʴ��duF�nRO|�v���uCdA��̎Hs#�EP���T�Y��m�|�YJ��6LLS��}PS�:ٹ����Y�vL�p0KE �ߤ�YM�/���K/VM!��,�S�c�9Ql�c����˗r Z�*���+L�9���NQ0��q���PON�%u�S�'��w���u5f3�������DC�;<*EC�� k��8�x>i_�~vy��-�f�@N�$ �vt��5�ZyMS�[��m�&�0�&5Z-�aHz�g7�#t���ĸ*�	f���М.���R����q��ˣ�^4A�➲�O,���>(l���X񟊡�z㴴���3Nv�!���s�H���<0�����i�k�嘡^��"iVz+4v�,�q��:re���W�P�P��O$��]Z>y󇇊�n^
b�ݢU&����t҃%����k����RY[dQ7GLp|}of���O)��|7*󫼧>�������VI7Zb{���js�L��L�g�a��Wقʧ|��\�>jr�=�Z��A'�ռP&�OZ�!��%�ץ�L-�����i�0:�1��l���TQ?y���_q���I���)��Y�^]�����Ks�k���8�8��_�I��8���-d�o0y���l%g{T�� jQtң"�W����� �	 �* �ͯ|:K�m�t�6˲aw��OrS�Wa��>�M�Cfx�)H
�.OU �f��S	��:�bQ����~ �%�i���+�0;4%s4��F�x�}@����҄����7�,|b�@��
P���~�9S�i٢��:eM� y�q��$�@	�xZ'� �S�QS��88�W3�w�;�(7��	��7�<��:+a�����?��!��>S�����`��f+?��8�Hb��oե�~��O���3��C��۲����QE��k9��K𔗤����(�
m8Y�����d�t.���\V��/���+���GΡ.?�J��ioD!OB�/"�h��9�#L�Vm�t�+���������3b��_Y�<Ɣ�a|.Y$S	Ŵ�������]�_��萓���NG�����<��A��<����"�bP��Q�+�5��[���yē9v�(�J����Ls������o����:�WU�z��Z���Mm�����Ye3У��P���Yo@Q�q-m�	��:ɳM�?��P��lM��Q��7�� +.�s�M@ ����*��=*{�+��!w`Ox�A*&g����q9�O�!p@K�C����B�K����=�V�)m�������)�V���2���r�j1ѡ"�c *�2*�����4�N�l�44�{2Ŝ26K���?/�CǼ }��w��C�obոʃL
DAMZ;Ȃ�}(k���"E�vi��M�.�y��U��ռ�Ul;�<(F�.Fy�=���d��P�!���+�`1�r�Ǔ��&�jhn��<?�~�IEg�?b�@%Wy�}*�_8U.wI����֞�k@�7��a"����΀�,Rl�%0�k�]�yDd��2y���Ům�^U���eB���V���S�9�^ɒ�x0�۪>�"ޏo�}a1$���ģQ�C�ee�Z% ���3[�-g%�i��@U!u�KtŁ!��"����Iձk���TU̸��|//��"^-D�uHH[6�y���؆n��/B�1��ȴ�B��$�̿�	Q�q@���Ǻ�E���L�����È�t� ��І��x�=W/[uIǛ����q��G��e:�X^J�����PXB�8_'�]�AZ[ع�'~/y���Z���K)Y�ٖN�	�S/��cNÿ/��ѭ!%̣Hk�^X_K�J]`���&�R���i1*=� ���{�Y�l
�A/M��hޛ��>�8O��!I���CP�:���^�/vAI���遆yb�=���u��nC:������h���$Js�	J�KM�#�(�"��랔NQr�1��	q�:�,�74��@�w=�ބ~��0wY���܎�vˡU҂�j>Ldl��w և[g� ���A�a� æQn�����_"V��C�!��t�/�h�"4r���wQ;3W�W�sCFw�I���#�w%�:��_+"�v��e�$��$�q��p�6GSQ����Z�:�>�xa����V�������:����b�`�6<��3�����+�����H"��G��&?8	�x&�a�+<H,ؼ��B����D�mH���
�����{�i����H�4����Z0="��1�4U�[���L������5���_n�����&�?j�:u�4�+�Ь�e=u�{jc�d���4G˛�᫹!�"��eӨ�'\��n�2<�2*<&���_�N��K/�����0ă���b�y��%Eulՙ]#ɼ�J5e�G��UuE�_X��?vm4�׀sA��t������ܕ|L2=h���Cwq87�a֭Ƣ�����압Q>�q)ފ&ҥ�n�L�-G��я�SI�h|�$qS�F�p����FX��:��ҳ��*QE�e6��߸h��6��;�I���<U�0�Q�=4 %�D����,�"
��F��g�>�I�ʻ^�q^���n��xQ֎�XoL��HSb���,�t:#w,{��r����Z�.��$2��ܟ�XS�ǰ�%�T�.o7�$���ozy�٫Ǒ�n���2S���
���2ҹM��ql���<z�0`O?|rDP�N�+{���b�L�"�pJ�����lX�����<�xh�DzzM�^���-x�����Q"��ztk}�����v�p�M1Tl=���#���vlp���G}�`�	+'�^/��!.$Y��<��@�ϼ1�{���PRԋ�_�{�yC��@����q.N�کM���ω�"h�;>~���s�|�&4��ݴ��^�{DO�O��-� X"!ˎ�1P}3��"{K 8}���kC��gw���E{���޺"G_�!=�������Ǜ�-���M�s_�|���n]�w�4��m�;<<��a�"�(�F�H��G���+eG��J�$�؀��v��"~�#�_d�u�e�1���B������IB�� �~w��pbF�/�
xk���o��;����$�d�
��/s�����ӻ��#����w�#�(:�3�R�d�oL�r�0�l]'E�`���J�Ru������3볈�q��L�*K���h"=��p5th�{C�ԩI~���QN�\��m<�t�>������薋�]��E�����-���CY�����@�u&�Z�j���x�!�!D��y`&�o-���ɽC?�t���͖nhs.NP9���m�C�ի2�&G��J���t��<#\\���LZQ&�����]��S��(�΋�����y��5Ŷó�{%�|ބg��&c�I��K37�1ߴ }��x�9i��=L��3�9�k���g׀F͝�f,��>0�㨝��?����{�%+9Ԁ#92�s=Ḽ@�x4�������g�bZg풦�f�S 	j���Yd�7$��۱�"���"H}��vo����
Y)�}�/�(��q���$�;�������K̦��'��G��%��t���:����I7�~̨�w'M��'�;p��q��J��Z�2w;��q%�2���ǽ�P�:h����15)�U��ˌ���,w!�c���*av�C���Y �CD�q�7s���X����~|X@kq����B�d�~�Ws�X֘@x��kV�E��dĕ�Z���gq���qD�5/����'���&�wI�׍P��ȍqFr �,��>B��lS�s�m�}�V0�.�F�T�l�!�i�����ީ�S�O̠��-ۆi�+�}PƘt���ܱ_��$���m�?E[�%&i>؅5}ɎP� ��Njn��r%~r �t�f9i�I������z�n����#�cč��,���C��f;�M�r턶�'�C�}��vn<qYR2�=os���vT�Y��.8�R<l�b@��F.UC�W�`�c`�W��X���Z�0	��x��P��ᾈ��u��A����d��y����.�`n��H�m_)&;�������|=���c����7�g�ix`y�)Y�e/&fBddi��K��	a��T�$�,���P��Q-��l����A��\n�9���p���*��X#T��C%����	������F{�O�4Y��=�
y�u�P�k��%���@�AN����f�	mE-�t�T�%�=���j�� ���(�i~�	�Mi����ͥ�J� >OSp yn�pH���u�,~c����p�O��e�0)Ȭ���7yex�/u&�5����-��xk�Ғ�R�8��J�4G왵�d��E>^k#���^�2FWڵ���[���jW��#�@ ���2^!���S��cF�:�>d�d �9 `p�w��b�<��/��um�~<.L �`�9��������|�_q3�%W���ri3�[Y��,�d��e���&�d����H��aD�ex�b�ұg��j��Y���׃�Ijn�[3�T̢Ztw�� PXqyb�9
��;Β<�"I�j�6!zB'n��a}�h?
��^.��X���<���`T.�jw0��$8��6O�l׾��ƉѬ��Y�``Z�D� �I������S�i8� ���7���á��Fת���Z:x�����B�fY�,�:�z�t�Q���,\2�F^:���ʼ}�&D��p0�Mu-X�.�����'I�>��)/툦�t8�b��b}ǟql��l�etA �X��O�E�%��,OP<�R�S[]x������#���k8�	��>@E|E~�
���E��\�]-��ί~��}�=tK��$�˕վoD2��Q�r��2�%�E������ݕ}LEј��Mb�h;�P
HWy]/Yd��}�QS�u� ���r`&)�,��Q�	��8�t�jξ�x�),COyI�:���xe���A�Y�K��j��b=�I�E�^���^0� ��$��>�������n	�Of����7����_���� �7�/���-��VC�F۬�u��^���tg�i�up����ɮɓ�κX�_�'�[��h�A:�ꏅ�N@dOY{;W�`8����MrJ��VI�L��V�o��v�Q�A�vљ�;(�o�a�6�&v �"6hfa P�b�]P��`X[�0o��dQ��tk�M,�n�fn���Z�`e����|��I��W��>��>�K���g�?A�0�I�6]"�S����BVgp\��/���&�
�W쁮3�cFe(��oR΃?*
�,��O���:>͆ 6��'�)H��nxG�c̎����&b�3P�ʧ�����hC��գK�[P���	aD��'^h��TP�^����8l���m��*~nq���L1�%+�[w�)��*�l�Ha2J64y��޸�~�"��Y�Lh�q�a=2����SyU:���'6�tUpN�ڞ������D��lxG��R�����DS��z�g!�Z�tV��T3���d�N��x�L��� �_dܡ�~rx 0��M�ۥ��b]5�������]��w��%�%0B6�Oi�U���%"�>?|�۪8�iT�7m:���i6d��F�ޜ����RѠ�e�O�}�lɺٟY.Ns�=���'dQ�l��b`<�37���D���a �6�A���HLE����H�#�Q��H�@]r�$9���n� H���w|B!�-|�+r�x��?"�j��o��M����5�F��y��T�����Xl)���0��4�x�R;r�F�jU�?��җ����>� O�M��=[�O����u!8����������vG�O�󤥚Lq�4��'G]���PR��H���5�J�6)Kge����3�SJ��vP��&˪�͘���Q��{��dhO?�t��ɥ���{U#g3�먡`����b� �X�k8����|}6�����&�Uf��(g��p��W{f�6�*%�4�;��?���L��`e_n�1.*"��#�l��61�GqR���۵��������s��?�v�����y%e�y�%u�dߜ�U�7R� �		��-��#� ?ͽ����l3���a�0����;�*��,�v��駓u:�&�G�G�<�9%0N,�ǉ#y\�E�G�|:@��e	��}�ϰ��DKX��M�:@q�2�k��RPH,b��YiN�<&K��C�{?�hGƤ�?z�ҟ	�a��YN3�g)�-�J1)�����1Xψ/��oi��s�CdH�vn�R�h�<h���3��
�IJ*}��eʒ��n�=�~����-�%��f=�����䒕1c���Sh�l>R��*-�sq��	&�μ!�͞1���`s�"e*�Ӯ�>��Ǳ�*,���J�2I�b��\�f�~ѳ�Ϩ qޗ�S�u[�ώ�%#Ժ7�4���o��[��Af��Gg�}�j8y�WD��q����83+c��.F:�Z�lH��N�3���u
�~�����7�p4	�Z�g�$�����s�&6.�2JA7�G}s.�B����7o_r��Iۧm��^:s�ࠂn&�D֐�����~Gt�F��z����8�uh��z��%�>���-�{���=i�N�,�uG�Hp�$~�C�Rz�¡g�N${�AH��/K3/=�x�.�$���3Z0�}�f!6��>_��j�����M$o=P��B)��(`�m�XjJ��\�F�ӦN����Cpf~����𲰟�S��V�6����������g�M�φ0�Lw�� �ިZq��4a:�P~�e?H�3����?	P.	���4��"�ӣ��PJ��V�N���KGnóS���Qkn ���"���#�cj~��^C�������l��<5b���r�x�>ѣ�X�s�ra��܌aar�؆论��hy����X��M����t�M�:�~�"x�w���P�Q��Pna��	j�i*9cx������8P�l�̳	%$�o�1fr39D�ň�?0^{���Zv<��j��X�ذf �eC�)�i`P7�V9hܚWW%v)�5���E�Pv`Y��5f�ћ�:�c˝�'?P�k�H�ge�S�i��<3��'�FJ�|�}	a��.��h�V.D� ߢ&W�>��UH[���Q{���13�? Z��8]���5,;�;Y�e�~��Vr$*Z%@6�=^��&�JEW`����R>�4̐=�#��)W���@��MCjYJ\�!�)��{tE��m�o��w�*U�K���&8c�HfS����1��jq�,�wK���.�̫�wî����m�L2�_a��L ?v�ָI�Q�=|��b�g�"����h�¥� ��+�;Z1,���r1�'-X�j�w߄���<0� ��a�|�nnJ���LS}�ot�݇��F�	��xxȢ�C��og��85i]��Z{L�eV�FT�91tۛ@�E��Tۖ�Vh�;w�!El1QW�U�\NyR>�Z�>�m���ԇ�yq`� �'	z(�	�?�]Ms��ήߑ�![�FX�:����t�ٰ���ڻ��F܌��Kt������z�Ȝ�,+Ԍ�"��
J�D9�3�>Ű��-��I߮F��;6C��Z�Q�5�|�C��y���o��i�ƌ�B���U�����\�I�RZQ����~�.I�ӏ��X�F0�$�S���_�H�Q~������Q�{���|��{�_�\z�;���AG��v�����~dk���y܃��'�Va��x|Hb�� ���6bp:�:���?��A0���.��J�s�] u6w.�	fӳ-���t�EC~��Kش�?5��-�B
S� y-Flu;(
P6�ucT��'{��;��B)B~���$s�, �v$?��k)�ޘ�\�z�e3��\ăl
zG����]��zI�2�7M�v�o�sT�y<����%᭄�֢C��I��q�t{I!a����۹���3:]e��-�I�w9e�����s>��t{���b�B���4����Cy�}@9�bDg���Wc{�R{	\���>��;�h)1�ڞ��,[Ϝ��|I�2����>`W�>�B���L���m��M+HtÛ�t��^�pa1��<���FP�X��-�L!V'�oK/�{�r_�ա(��+���Æ$���C.O��|��MY���������GFlQ�ʩ4|�&�a�+�2�e��B�qY�!T�%r�-ўo�����GJVP��a�ut�B״��Mt����x�x���}��^䱈��J�ĺK.K�0���j.ڪĎe���E��KC;�(�fm%�AO���eĕ��.�k`�^1�ei]���8�H�x��N�#���Ո��������lbn8������.�Q���&+Yĵ������#��G�6�&̾�ƿ�^��i;"�ZZ����&�pj6�aG���rB�<���U��Rw__P>Qx��
�
r�Q�?ʴ�̎�]��I�.�GSiΚ�3��B%�sݷ>L�}�Jj�8���p_j�ӂ���0�f<W�F0�F�r�{Փi��C�)=��Όʘ�����KC���#�~��U��%Qu��i:���Q�~�&�y~	��Ϟ��E��;;�3E��	s%-��[|�1肂N�S��o�t����z�7�U��p�ۂ���ʨ�$����m00<�j�~��}�{l�k}- 6
W�2�7�7%�C�e��O�&G�g}�®���UE/V6X�wxvU�ՙo6���5����C)�~ C��,��N��(�o������_��x������:�u�<[Ur��FA?���:I�#��
�;_l�+,R��.m���`���)_�Ȉ��g4���DWc��ۉ�Wi�6��ḟ�=��o��+2�_�Ju�t�ag~�"))�/Z|�m�	xMPM?E&[�0Bs���E��_z��2���ԧ����61t�]�+�U!�]��rd����b`�)�_k4`?����z�_�r���=L沢���sTX�I�\���x�����y��`�_{s�z!��h���F٦��I'����d�Τ=h`���8.:`7�tgo( �A3�PX*����x�×��|�����U}s[��4���KHx&�ُk�Z�pd�����z�����ӻn���*����b���f��en2�:R��״��쁔gi@�Ҡ^4dA�L�l�2�� ?TB�����W�1���>���|Р3IE�k��
�N �3BR ���;�q};�O��	0+��0US�Zה��S�h���f%����/�Ql�P�?���s:*�}��A�ck�R�bΑ�g)���=��	�U)�΋Pj����:�k�*3���dl�
MF�T_36�n���j�H���-_�p����)9a��gH�1u�Hq$��`�t�֭
:
D�C�V��&�Di�@������h���Z�(\Fѥ��0�l9U�c��>�u{n��,�h�p����c�g��i�<�7�f��PEm� �xp�ij�ӛ�5��C���M�1AU>�o��w����}n�?#Ŀ�(�`�"]�B��(9�X�g���b�F2T����7�r�����8�K�K� �%w�#k�Iv�;n���xC�w�ܟ@�O-��iĲsAW9��W���gl�t���h��^�c��|"��;�xt7��Mc�C��\Y����
i׺:G}�c7F,�DZ���t�x��0RG��	}�B#ٯ�j�Lq�^�������2��`+�#\ni��ͤ}��3�6��RD�$�2��� r�Ե�O'�;]�'a�.9I���ϼ �3�Ȥ�񈭟���-����<@F���P���m%��V����̩��'�Fn�*ݓ)�E�j/��A>�_�a*G�A�|�f8�m�&>CZh(4��k4)���i�eI���4K��ȫ?�y/���Uj��=�yxa�|n9y����/X��0���-'x"��$�����.���eơ��~Q�Ѳ�_[9�7�]ƪ�4�]h�=1��	��x���p�+^�$?�?8����<�R6�魛/�$$c�CF?����0w���N".�A_�_�����Dm�cFI�w��t�(zuO��.
YkE�k7��Y���aO>-����9>I���Mh��P�v�O#r�o��T�����������!�D[�%����%���:?CgD�a
�:��Y�T���
a�G�V%�>Y��*�ȓ6�!�X}!=�*�Z	�!	z����%ƌ�UO`�|����DH��$�i�CB��`��`B5�y]�b�q�|p�lĖ'=��D����_Z���1�^�?7��7�R��0�)]�����))%9C%{)�̖��gK�}����W�f �X��(cME9�&!�}�:l���F�c���pc�V����,�p�
�N[����{�6���gE���`�wѱ�f��a{���~�>��@ɝ���ՠj�^"͗���I6�:ot�M�f+��#�!����CzP��3�RɑA�'6ޫG<7݊Zm���8�"}�ܹd��)�BJ���tO�i Ɖ�#0�6L��V�x��C��I֪V�j{]�0�W���/�uG��������\Bz�EI&�І�@%���DM�U���\u�$G�fxm��6j���{��ϞOR��g��&X-G���$ŸX�@���K��8�VL�E����}�71*�}C-P9��"�hr�#c�P�g���8���RQ��D�8 ��f��iz�};��7L��;ߝ��\&I��_E�̺6���d�^�"��e0tٜ`�ԊոT�~LRt�'@H�&�M�T�Q+͜ ǟ�p������x/��0�dz�I$eܤ�X/�~�S�IPX	�����>Q���$�.?|����mS,w������R q'�؀���K�X�~;�|�b��6Ö�
t�f7��P�펧���Ƈ�7\��(�Z�+$���iL���~+.{f:C�#��TK��h��.<�¿ ���@����&�-k����KkȾR26Q�XF^��oy�׍J\��~r(���J �k��-�=����	u*���l��� �Ru�BeS:v�Y����:�����¯��Q9�$��|KvDw�4�gV���F,6��~^M�_� �jM��v7qd����|	�IP����� l�NƉ:�¸;�}��v�+��� ���J�"3�:��dgc�|�t��BY��+��֬S���oT� ce"l�*�+����*�v���k���8A�@�j�K�Z�-�����>��]������	l�W�O���|�\�r�)d�%eo�������^i���+bؓ���<�;BS�A>o�'�!��p���ՅG�:�f�>�7UDӇX7�&�!�q�B]"�q��$��M؄N�����:ޭ�?�4��`3�F�-�HܭZ���y�C�^u��}I�`���y��rH�FC6l��P?����ʆ+"*��D����/k^9�;;c���	��F�Ĉ[�܂�
�O���Ic�7�-�=�e�6l�U�Ω=�;��T�)��J� �����y-���A�8fXl0�����K���G����P�ܤ
���LN��*���	$?Ė\�A5��K�����                                                                               
     �               X  �0  �               	  H   p�  i           P K F P Q S N F       w�Ա\���ݓu����3c�q���[E����kb|���P�>�팣 �@4��,Fȡ~��2Ɂ��Ya~y[��Kā*�����햢��n�4��֩$�AZ-���d�������W.B#�ݧ��¾b��}H�	�D�.]��1k�,K#�>Rr�? ���kt<ӳ��F�^EQ)��Dl}@�F˘�G�9k��Q �&c9��.>KPA��j;���da4��<��K�?�'��VL�����b��ےQ2�N��c���,\�m�ʝ^H�y��Q}.�8J�ڎ9�UN���:B�l"'.�?7�	�A�}�dýL�ǐ����k�/�u����N��>G���i\ ��|#���m�hͰ���yU>�4�a8#c�sj�@����>�QDt,5#;�_6L�I��2�Y���Zvd�8�8�Z�H�_K�����!u�bu���f^1=�7�%��-z��"�f��b�)�W* ���.h��]aw�ekdq�8� I������w[:����$.m<��Cu�~�d�n��a��HkƖd��G�'���~t�yV=aA��#V�K@��qBb�`����R)��;�{�+�Z�xV��,��}@ٞ�j��?��|<A�e^Y����q��u[��{G�ތ�SϴK�(�	�Z�P6�-FR��q����(����e+ź��=�{ٰ��`vC���;x��9��_�|��7KB����!2g��g��AF��]�h���C�K�Γ��UA����A6爄M�c�d%nQ	#1��.�ɺ�ȏR���)V=���"{z�ȍ&Jcm�b��?z�+/����U���e�V��C2���s������Z~�/ك�^�	��fղi/�u�(M�CP9z{̨~s[�"Br���~����u�f݅��x=��N�h 0��U�e�-kg��`��ۑ{��UHt>��K�n+�W�A�n��S�&R�5v�Z��E�V���.��({؄�Bݳ����Y��P�s{?��������x-¾�7��9rh��g����K�`0�	J�AZi�
����H\���R�>��:���b@G�Ɖ�*�Q����kj<�L�y�2��r��R���                                                                                                                                                                                                                                                                                                       (�          d�  (�                      q�  ��  ��  ��  ��  ��  ��  ��  ��  �  .�  G�  Y�  g�      kernel32.dll !FindFirstFileExW W CompareStringW �GlobalHandle _GetTempPathA <FindVolumeClose �SetConsoleCursor �GetWindowsDirectoryA ^GetCPInfoExA GetPrivateProfileIntW 9TermsrvAppInstallMode sGetCompressedFileSizeA   GetCommandLineA   ExitProcess   GetStartupInfoA                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �W[YZ[X]^_��bc�efghijk,mnopqrstuvwxyz{|}~����������������@�����,��-�V�%��m����ֆ����������������Ҙ��՜�П���㩪���������������������������������������������������������� 	
 !"#t`&'d(.+�g01234567�987<6?@IBCDWFGHIJK�WNOPARST5VWXYZK\M^_`cbc`efghijkhmnopqrst�vwx}z{|}~�������������������������������������u�������m��󴲳���������������������������������������������������������������������������� 	
2i{gT!"# c&'(9*+,;./0523456789:;<=>?`AB#j!'3)IJKNOP1RSTVWXCZ[\]^_`abcdefg(ij+Bqrstevwx�z{|{~�炃������������Б�Ӻ������������q�������Ū����������������{�������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRS�1r �=~��9z]�f�ptfggǒ�I�U�T|vw�yz{|}~�����������!���٢�p�������,Ƈ*(�hb��ծ��pr�\z���4ޟ�0ڛUL��Ɩ������@���\��X���1q���S���o��k���g��g���
{���w��:s�$���]�n/�j+��v7��3���z;X�F��B*&���3?/0�V�R�^>US��`�rc��HKL�*k�6w��2sZkox]kD�Gk�C��On��apq�P�\��X/N���@u˥>\g�������N����(������z���!Ɋ�=Ֆ9ђ�P����0ڛ�L��sH���B��$����\���X��gT���P��h���������a���}��y���s���p��!�f'�b#
\��j݆�<5�?0"���u�{'�G ٫C+��,./��>34�R~�^��ZB�&g��Bc��AKL�*k2�6w��2sZضS]]^��mbc�B)�N��	Jm�G��uuv�]m�Y��䥀�n����詑��q𱔘.@rǖ��ą�.��Q*̍��%��&��Z����:ܝ�6ؙ2���<t��������C���_��?[���2}���R�žn��@j����-#����Zy��p���� �����h)T�t5��p1�X�����D�@ǪL(.f�-x�6�{389�_�[d��'`G�lM�۳���4u&�0q��<}X��]_`n̛�!B�g�1����[|qr�Q%�]��Y|8h*������ ꫒�޷�}%igf�����x/ǀ�����C����=Ֆ�9ђh5ݞ��oW7���I��E��TA���]��/]���������R�ŭn��Uj�������}�֫y��]u���q���&�!�,-�����4�0�r3+�~?Ӑz;"����ګCL�O��K3�E��;895�Ĳz�N�"BEF��DJK�)jx�5v��1rU�S\]�;D"�@��Lk8�pIo[TB�p@Q�\Y�X����j`���
쭋詏����������[���ą�.��*̍�C�QQP�J<�.^���T����)��e����g2F��B��c�Q�(('1����S�Ĵo��Hk���b��g������{���w��s�$���0	��j+�v7����E�A��M)i�c(01�W�S�_?�[d��G`qFcI�fo������YST�2ss�>��:{b��def�^��clm�T9�P��\{�7Xy�����ࡑ
�a詌��n����q ������/ǀ+Ì��������\���4ޟ�0ڛ	L��������"$����~)_��[��I�^f��� ���h���d��`���r2�5	t���p����f'�b#�/�9*����q2q�}>��y:�E��!UG]O�.��нU7�Qɵ]9qճ����'`O�#l��/hO~du Uar	�aW[\�:{&�G��Cj>[WH29^DU-�����wׂ�Y-��3j�yyx`�����������됖������|-ņ��$�*��FEINM>Б�:ܝg6ؙ��������J��F��kB���;����U���Q��$m���n� ����`�ˤ|��Zx���
\�������@!��V�����%+�}>q�y:��E!��,)� ��ѢT�P��\8�X¶te�_`�*EHI�/h"�+t��7pW�Sα(Z\]�;D<�@��Lk9�hI_kTB�ppQ�\>�X����j^���
쭈詎����"U~񘙚���ąs.���/���C&���=Ֆ�9ђ5ݞ��oW����I���E��A��Ͷ��|<�+('T���P��Ql����' ����`�˵|��Ix����L)o�� �f''�b#ׄn/�B�����s<�8�{#-���R��֧O)�KϿW7788:�����%fj�!b��-nI|rkZnw�1r"�=~��9z]�/����C�O��
Kr�&w`�x����XE��K砇�u����x�jlk�8o�����o�'����ND���&ȉ�"ԕ&>Б��Q+����8N��p�Db���#h���]���Y��)U��ٌT������$���e�Τa��\}�������t�ߓp�ۓ�f'.Q��j+�v7�r3qw,��&�!�L�H	��T0ۋ567�]x�Y��%fA�	j_�[JKLB��v�[��_XY������E<� A��Mh�8Iz��{rs�RE�^��Z}���o�uut����������w6X]\)���%͎[!Ɋ��Y�HKJ;Ӝ�7ߘo3���O��9O��!����C���_��[��ۈR������0���k�̝g��cc�������z���v��"rd% k�j�%.: )=�=6�p1s�|=��x9���ܩA�M�I
-` 6l>2�].�Y��%fA������.oX�*k��6wVZ���R[\�:{T�G��Cjf�'xy�\rqr�Q!�]��Y|p6ն�l�{xw �U���{)ged���-ņ�)���� �����$��?א�;Ӝ7ߘ�V38>=N��J��cF���0���;���׏P�����T��o���k��`g�������~���z��'v���t�%&�	
�h)3�t5מp1������z;"�F$�B*֚7,-.�:�Q_�]��Y=������"c@�.o��*kR��wtTVW��R[\�:{�G��Cj���mn�Zsrs�Ru�^{�Z}�7PkQ{yx�������]~�`fe���ąZ.����!������Y���>Б�:ܝ)6ؙ�W�:=<I���E��1A���[��;�.)(U���Q��m���n�� ����`���|��x���q�������g @�c,��o(j�P!�p���|=H�x9��D ��-Ή��զH	�T�P4�D6�w<>?�%f�!b��-nI�z[�A����2s�>��:{bW#��<����H$�T��Pw�\}���������7
쭈���g�����������\I�Y[Z+Ì�'ψ!#˔���\@HG4ޟ�0ڛxL��Ɣ�r�g*��������fP�y�������3�.L$���-Y�f���n���������v�ٍrd%��`!oT�}��*$5�0�r3�~?�z;"��&$%�C=�OãK3�k4��189�_�[d��'`G�|]� ���@���p�Y��[Z[��__`�G�C��On�n#��gPF�|L]�XQ��W砇n�svu�����uqmacb���/ǀm+Ì�'ψQ'��8��\�BHG4ޟ�0ڛ[L���D;����#����]���Y��eU���Q��7����i���e��-a���!
	z�ݢv��Trd% R�"6-�(�j+a�v7��r3�`���{	�G ��C+�Oѧ#ټ��ʻS}�_��[dCÇHDFG������*k�6w��2sZ�>��B{aUF�PA�L7�H��Ts������]H�Y��䥀�z@������fg����������ɑ���򔲃�A8VSR#˔�?א(;Ӝ��c,L�6������0���G��C��Z_���>�"&%V���R��Kn���d(�>b�Ք~��jz���v�#�<+�)�/�-�#�!�'��^�����s<�8����������פN#�JüV6� ��::;�Y"�%f��!bE��n[MMN������1r4�=~��9z]5���bCYmNX�fjK�V1�R��^y��~��������I����JcL��JPZY*̍�&ȉ"ԕ�8��^�CFE6ؙ�2��N��į&�m�E�����Y��X��T��gP���	�k���g��c���u��x�Ӓt��dp��������c,"�o(ڃk4�G �����x9<�D®@$s�A++,�JC�V��R:Q����+d�Ng������.o/�*k��6wV�zs�=~w�9z��Fa������O�
K��Wv7������Y&��(ࡄ�`�zts ����9���`�$�+��.Z�!�8[�� ��5��8ғ�4ޟ0ڛ�)����K��G��WC���Y��X���T��0P���	�k�̊g��rc����� w���s�$ �g n���Ɋ8)@6f�?0AJ���{E�G ��C+h�	��нU'�Qٵ]9k�"Auf�pa�#lB�/h��+tS�n����<}2�8y��E`5UQB9c]N�Il�Ur�Qt������Zm�s	ᢅ9�����x�glk���� ���ɚX��-m*��B��(���3��b�^�� .Q���؆M��D��Х@l/�[��^���W ]��۬ll���'���f�Ɂb��a~�������q�ڸ�e&��a"��.#������\=��>����^#$%�CD�O��K3f�>��ȵ]�Y��%fA��F'HI�E����4uv�0q��<}X�YJ�,����B#�N��	Jm�5v{�����_+�[+槆z��a�ssr����
�[�u�q_^/ǀ�+Ì'ψ�%�����]�XGF7ߘ�3��O���K��!o<32C���_��8[��۲��^��=�Z�g��C9�*a���{��<w���}?�����c,�o(�k4z���"�=8�
;�E�A�M)����ϼVF�R��^>h�d@^g�qb�,mQ�(i��4uP������=~O�9z��Fao��Yhij�I�U��Qt�������V�������>�����D��x�elk���J����ԟL�[XW�S!Ɋ�=Ֆb�0KGFRJLBA2���N��J��ȭG�&M(.-^��Z��dV���R��j�����n��a�ʾ}��By����p���f'�b#
��s�t5�p1��|=�9�T��ݮ@�L��H	,�TξPʾ��Tc����ng�9���N�xi�+td�7p��3|[���E� A��Mhd�yl�g���tuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRS�v���T)����1qC�$?sܩ%F��o��4��v9�ܹ\_'�z����� A�h���ƫF�b����;4�+�C���+�`�RJ���������C��$9F�o�3�h����z
�"��f��i\����B\M�s�G�>��}E9�j�]�^V���Y� ��O�@�Չ1�qY?K��֕���nv���iu��6�t���d�R�_^�U.��@e�p�z��m^�#7�� !�O�V$��e�@��|ykq����^܌��\.C
v��t�T��'��mu���8�k;9�SA~!��!�M���0W;�Ӱױ�t��{&���<��R{�}Q�M��;��*w͐P@%�Q��s6 �������hH�Zx�m��*�@r�8��D3]��(kU�to/�uyLUzy���z�*�P��ٯ*8��<U��a���\Qf����=֔��ö́�M ��P=�IT�C�vB-x2��rp;>���x>y�]~5q}0����.s�:	�/���}r���N�L�n]����8֣���F�![)v������
S��B���L�9�Ԍ�AZ:D����a�?Ad�;ƶ:ƴe�7;�5�%E댛c!�ܥq���E5oE�h�ܨ��K�c�	*X+O��&���G��(��і�B:O����4Vy��r��Se�����M�yyN'�y�l��հY���jkO ����A�šR�S�j}�[U����#��÷s��b����Wz�d��3�Ž����x�"�u[��aAn2���������b�������Ꙭ�A��'�D~�Z*U��ԩ���&�����Ys��>\l:l�O��eW��l�U�4� �3ʝ�)7�Vu�>���(�*�5\M��-�8M���!s�<nZ_����|ݩ�nj���|�C s$�7�m�_�$�X�(ޏ��*/��j-��Qs���:��b��d�~u�-�'��ͳq�5�a3ẶT1�YO>:9�y Iʟ�^����ӌoRčL ;mTOmc�>%�M���Y�@cR�gӽ��Y�WxS�N̝��[��C�$o��ͰcQ@_@���E?d��� �a��"����vd�͜%M$�;�TO�eM���Q�B�^���}ThW�J�8��=����+�h��,x �X9+틜��2�7�(I��y=>|�_y��!���`��~�&ίB�W�=�.�Hc���T+"I�8�[QcR��hB`8e>8�(��;��_ꜰ���}���N�1�Zӂ�H5���N&,5�tҮ8L�!:�BR��5�*��u�;2�#��h˽�J+�:��K�<�H9�L������zC&&���#���!]���A�N`�v�Z �2B��qm�������'W�oM;��Z�FǼFW���&�J,4�`wFi�	=^:-�O��#T��� ��ndX���iҐ��45��5s����g���%�tf�R t}X���S����33p����������i�O{j�Vt8���7��	���Gcf9'���e�f�ͪ?JJ�Ŏ���ֽ�ƌ���;Q�鞴�[v�\m1Ꟶ�g˅���x����D���>�D�� i��S�t�՞���Zgm��{��wp�I��"c)�U�4З]�ɟ�cſb �HP�^����wn�D[�yd�@/L��D����������,x�M�r^�
\m���j>_h�ܽP΂ިc��Q$_��\լa���.�%������]��2�qQ��^��d#P1X?&Wm���	F'2ԚߞZ&�5�7)�j�$�]�f0��1L�Qu�ZV�1�R"�k�4-��<�j���ۛ�SU
c����N9�r\C�0q%T[b��	�������D��t��c!�W���� �`�D�s`+��.Rq �i�"�Y�3d�^�A�����(���]T���on��
N��p���[�]Yo&�6�z -?DSA�m��PY�բ%�r��FiIm���(/�R�E�ǉ��K�J�]�ƄķO!hk����ln������e7I1:�T�H�)q:$�h��ͯ�G��Μ��U�{�p$BB�E��*�C��ب���Im+<f��/��G�Qm���K��bϷv��r�i/�2��ʠ�O�e���ԱY�=�,��j��ó�����F</)�+����7'��[<�Bpm�ڽ�&���l�Kr�~�w���Y8F7�q��^8��i9;ذ�.7���D�@�"u�<`������c\ƹ5Џ!$4�.��T�f���[���br.`��DP���0�Ε-M���j�B۱�8�6����$Mb�����,��2���](���#z�׽s���eН���Tt��)s���N\�&"��R�J �jd����V|���T��֍�C^�8T��^�aT�����&:SwBPR�sų-VD)ф1h�jK%���%�r��&��||��]�=�K�蟲.�������N=�k:��;�zM\����+�� t ��,X��+N�t�K̎8Rⶎ�����`dk�Ǣ�)���@��ʵNE��04��-^��
׼*-��`E'/<��;;�Y��*����n�yX���G�ps*X}&���m�4��/!��˛L����.h�1-��6XR��2���Ц���/?S�,x'�i�G�K~�e�G��[�=w��0R�J�'��*j�1����_�d`�M��I4��?<e��Zx��&�M�~�'���${%����"o���	����0�o�t���lˍ�\�����,����^eLC�c��_W �٢D��3�~��āK��L�!�9��6$(�~).��BF�t-�x�G���m
o��0b�)n���q���Xŧ�	l���q+D�b� xn?i d>nIp�V��*�>[�Hlh�����E�@j�&�\LY6ɴY�1�_��[�=�E�R����7IL9��i���Қ����T��P�M����/�K�2�(�%H|{V�}�A��J�����u���P���
!�k�{~;��JҼ�#�/�G��U�F�������|zU�����1�cS���{~��"�@�p��,2�2g��̑.�Aw	�Q��>����	�3��eї\C��p~|�'=�B�ր��YxJ,3�J���N\k��������C���� {#��J�h.����}�P�/5��5�HiP4�[Dژ.DJ�ź��]�`���p��T' TX�Q�X1R  ���뒲�9Kdxrh/_���WQ��a�)	������t:Oޓ����&����~�f����5@t���p���'���q�Z�V�پ c$`B
˟����.MmHBG���=F����Ƥ�Y�z���[w}�NJ^�ש����`.�5�!�pi�䧷G��ɜ_K�Fُ�	�0U�p���@�v�W�'���6���\2O{W�Pz�2��cl,J�͠͞�a]����,�^�_��V��B�?�t�Y�X:�0e�g^�3�zK����t��~��l�%����hCx	X��ٝ~.[�k��'���  W8Y�����)���'�#���~��n ���bL�Q:����[�0C7�W�T�9o(��m8�ө�5�LSr�)���;���Zs+%����;k*G�[>Jf��οy�V���}0+&5��x���NH~6g��OQ�g.!�N�c�\[(U�Z�;�hL"��6��Z	�@h�h�W���X�@���CO6�΃����	�z�!�/�Cdf�/.{c)x�MnZ��%,<ؕ& \��y��ਏ��+2��%�~��P��1�Զ��+T�t6�l�[ˮ�*�`��;/j�N�gh�	r=��Arbꉊf�n	Xb�6��
(c,>c�&LX���J������^C9xuv��D�&�;O��!��p��:@��I������=��^�%nO����8�d��q&�F�?`)Rk�;#]��bL	`���^���".i�z?V�����Te�*��ub�_̒f^�i�sW��uhG&�0��P�s��tH�?W?����0�� }=�"�7�o�����y�G-d���E��p �#��������}~��'c��~�
#�^!?kKusǄ��C[2a��X~�&}�{�*.���v =_@���|��]yN�5QSn;�t ~C���@�E=�f?�Wr�0�Ғ��GH�]qpw�NZ���`ޫ���}�"#g�p����f�e��X���J�;}a3]��k�Q����,�6��u��s�b�(ж>X����e)C��]������LV������M\������紝)�p���}@GDT�*$*u��z�>ģ+���� �B��BnI�5|��B�r�ӥ������R�L^f�l�`Dbp4hlL�j�O��	��I���J� �]\F�b��n&6��u��f 鄖�����J�M��فɯ7���t"�F� �q��ӡ�8"��bC��� �����h�\P�(8��}'$���.�-C��=�6bUo�Oü��8�/�F�/ٹa�/� �=C��b��D���2^~$�x�J3����y5�'�W��_�8?<|�d��k��<<nH栶VA��~;O���JjJK̜H���k��n]�u�g���/�h��N8�X�I5�c��^4������w�V���N�s��Y���*k�,��g��'o]gO�e��B?jV~@bUe=?��HX@ۆ�cI2&�p*e��g.XL��_��C�r#j�m"2�M��-�E�Ɓ��_���wR֩�K��=⹖����
MR����+�+m�Kx2��O�e�Za��\܊_�P�?��8���F�Z�m�1�*L������$�6H�2���`y��9O�+$�t�S��w	"Mg���ɖ�Q��3����;�x����@�h�`W�N�q<X@X���pU�L��w��L����E�}��]�~�y�\J�;����:��֓�lMi@��?ŰaJ8~EާNT�/)N���~S�ĝ��7�1�w�w����e���w�
���^��h�����%��Ķ�UgM0�	:���S��Yf��^ͽ'w��am��i���Ｚ�ꬭ�yC���P�v�fq�uf{�>�J�(��.b�}�%������YԖ*9�],W���x|D�L�Z9^"�g��I|XB���Fr�$��O����hzu2_���_����<��߈��$[�t,�W_Yt'w�S��H�M�u�@s���D�5ƪ�4&!�����
ɹ����ۯ�L=J�SL�7q��y�kHs���`6��sM��/(�R����&�Lj��$�*�]^X�V)�*w�1�+����{���l��8F���苀��7_��>g�������I�k�(�'�]�3Z`u���a҈,h��:��:<��D��^�m��^o#y������ O9Z��6��9drJgo{`M������0�8-� 
���Ԝv7���Bu�˴��0K����������:�Fq���<1z7zs\Ɨ'(�5I��-��R��F��g_������I�'�)%l(is��if��i��%8��?�
�M�e�W}��i�a~�u\Ɋ��Fc�@d��(�.�N���X���Pu7�*�2�'����RC�^��m>'������/3HZ���LD���ƭ�����$N��K�2k��^��M�nQ�M��j�I�cjF3�36_�e9>֞���a�,D�O��lb8�0�Z�rTO�mxK�s~���������p切S�M�K��M�&P6�����9�����CeO4h��Հ'N\��g�}�Ft��ZѤhBdؖ6̮{�� ;���D��L�XZ�S$ęN~4N��u?���@��K�ͨ;B�͡�����I�H�8Y��GB��.�X�Mv#��Pf�b���U6DC�r�	k�-�8^b&�b:�^4i(�(r�:c��mn:�@A��Zu�`�ȶV =N����<V�Q�}��]�^�8�����?r��pԘ����������&)?u�x��	�Zk~�=�wD�z�5��:�,�ӻK�)Х�q���>=Qh�U��2��D��q`�����Ջ��.�����QA�
�(�/f�g��3D�����9n��[��v%8�G%q�brM9]�5�a��ī$*�+�;fow�B�� O�h�b9� ��!���n�=�!~��A�/�����YX.~�dj	���&0w����a��S���k�a ������DD �� Pske��Ӂ&5[8�[>�f����o[rI(�0V��\�tb���%��7��T��5R�0�L�&gi�7��"Ȧ�?ED����z��Rl������ϪQ75�RJ��j�uH��8���f᧕a0i�Ě�Jj467
� X��%���$�tढ़|����:��a$A�$)OJt$z�2��,&m��'ƕ���"�[p��B��k����@��.�8'IJ~�l��w�V���<��j^�#Jr�]�,B���X1��R��s�y��f����)�3�{x�׎���9�%o�`����8���n��(�3��v���6� ���u8�*�����F��\�m����,�4yt!ϔm����Q�Ƥ��u�����VDE���P�EB�)�b�-�9�*2|��<W0[�bޚS����pۍo��^=k��is����B���7?q�h ���B1���
(�
�Y��M�Z��(t� |vT	E����Y��?�9Ο���k�M/�[��R�Y"��TK��I	HUih�	��,t�8&��kCMW�Ķ�:j��K�u�BK����d	��`kE�/�ՠX�.!ѱQO�0���:���|^K�V�|�c��#ۀyi�|QgI�R�sFށ_�r k�踣T��y^`f4����U`5�4��\��!|��tG����1
���R{��!{�_�X��Y��X�����ވ<� ��`�1?�Cݟp��k"Xp`⡒{;����.�N�}�z�{���<�WK����,�����"�WwW�������&BǷJ�Yh��u�:���H�����M��s��d�� �%?����(Z�9�R���7�{�l�ZI�2/5����I��$=awu[9Nz[�f�N�ls��m��a�8#�x(�KlS]e�-hC�EpZ�G�2T�e�B�C��s#=( �3���'�������mG��˫Qɣ q�E�m+�N5�m������ux����K��p�$�duO/�y1A�J,�;H��O��P��f��4?c@j,;4�ѿrbYu�Rz�F�2�KL��r�v{��� L��X���_L!b�_��}L%[<�K�!r���O������b��k�~
�6s�lPa�M��f�$
�F��ņ��>�5�E���?y���"�Z;9R}$2?BB�H�k���ը�-�Y۷%L��a�ȭghB�r͂�	�(|�X�r�_-�,F�N�2��NՌ����b�e���Բgn<�� h�o�\6<�t}&��#�}A5�AyP?M0��� �ABߍ���r�`S�#����[ې��Ay��W���w[W*�8Ƅ"c�C���z(m�1Ax��p��d�z�� A��cDJ�>g�0��[�狗0�~K���N?a�A,Ԇ�4��s���b����\ě��6&L%���0`��(h�7V��6�k�m�D��<��p}Dx@���E�fU�{ފ���V$y�6�SI/�.�>�{�:����]�O6�; ]N.�b���5b�Ě.]��(KXN�@��ָ�nF��_9�D�c�� �Co9�q�{�L�KJ& ziDUtc��Ǩ��M���� g	��zC܅N�6�C�����
��΃��YqR7� 14Hy^%t���Kp��yKo4��|��L�$���\$B����_7�48��(�$}h)Bj�����p��\���ڴ��f����~9��[�s�.�Au3,�W�G誥fZ)�D�����N��4q�[�vn��ZeVv��c�yH��
D�y-^K�mZS��>1{dA�u�����.��\�z�g#�*�i�뛟���8<?��<b�o�)D2Pٿ�t]�?�kr2�_�� �rQ�L���d��0�8?��M�a�A�d[��Z!��,�<\����+��t����֞jj��E�]�^����t_؝h�@�
'_	��|,O�)��m�N�25Almk'|2I�`��gȜ"ܘ��Zb!�0��Q߇}&K���'���
������ F8�MX�!낍P��#�'�e�2��2�#���ɧ����޶4�z�+����&.̤��b��^�< M�y�V�k���MY�v���a4�+
g�*R���-k���	#���Ba�$=�����r�^W�f2�2�OؖV��������j�_���BY�������Zb�լ$�ںD
�3*3j��q�qه���u7ޱe���/u�$���jf�д��EQ��}�W@�3q��v,#)�o�.(.i|?1��Rض5S&W�\�uvŋH�.�	�Uj1�W��t]�m�gc'$*�N�Y�����J�x�2�����~N"~��`WS���^��H��&��҄ҫ����&�OW�<T�KI�=C�^�̹�'�c?>G�^���y��W�TzǊ!�e8���Z&T$#ȏh��>KI~a��Q��N�6��O�0�vM�[<��τ
n�є�{�^�e�K�7�>Kg�Ht�:�u�$���k$Wn�[>�����{������1�U�=�ܑ'�C���Y�:�Ih��R�BdA���@��t��hJ"�!�V�sv�rp�11�YP��7���O�(��L��һ�0�㋈p��#Ң".��ϲ�6`�f����&)�b��zH�}z'_�2���;�L�
!����*��')�^��?6n���sl����T����vZ;�yb�>W*������N7�����Z$����viRo�����7b~
`t�u���s��E�e��q���
O��d�4��O9��*����������<Yg�8`?���8�W�j���F�n��

u�|P�/�
ǽֺ��O��@���ʍp�8�5źp�XEk1n��=q� /��}Y�I'��)�_�q����9 _Z����_T(v2���Z�*�LЅ�KY��4'���%��p�\����JU;��[$�<:GU�����5ф����Bɗ����#SH;Kq3(�1�\�s�����4&��iP ��\�|�X�-qN�c�0Jd���o�?�N ų��+�Ƙ2��k���\�s���S�� q*���^�`��q$���b�җ�X�j0���U	&�n��~�6ŀ[�4�9����[�U��'��:�����'��̵8��]�.Lq}5�X����#t�@W%N�RpϔkRw�f��Bs��ԫb�&�(�:��艌$o�h�!�:측"Gׅ��U�k96A�v
$ �¦zD��hA]�=pũXė��T�
y��	i)K��ez�Ы8�p���<9��-���|�|_q���rI��ƒ�
1�A�j�3#��R��V�T�?z�����Bӌ,�jO>U�Ò���?� ��YݶcZ+�qw,���9AO�R�!�޵�Ag��	�/��۾�|�"u"�|��Vz�F`U��^��Ӹ��k���E���>�9���:�g����U�a�@����Z+��z"o)�ݕ�f��j�ǜ]o��l�A�O�����`��=�`|���-q,���J�&W>AF�L��[�t��X�5߰͏C��s�Wo+R{{P�w��lWA�+f�]Αxi�V�]�}?xҷR����$��6��?<�&�v�ğe�뭌�|��A��Zξ��|���TT���F�eé{C�9�Q���xq���O�kK��Xkv�^U�S֓�H�'	;������<�TvGd6_�?p»�d>�ٿ5J����y�Ϝ4J)���	{F�TA�[���=3� ����c�V�b��]t�B>{���R�'���Qx��hl��H����.��T��:�0�����o).��8�g9?�0������r������C�L'0+n�]�NAOP71�{3�n�.��M�D�ɪAVjGhEQ��e~tY���M[lY�{��B&�
��g�������P=��}�]�Hs�)y�<I��=�6z��$٥�k�̵/m�L8�Z��Tʚ��|X$���/�O0���VtB3Ka��䇸\�%�)������?�W��&�R��GSV�����w���S��r���:��	���?����m�׉�ϑ��K�	;)�T�2��.�P�h\�i��5�g�r�z���!B��Gg�,Zq�s(�#�H<�X��Y�]��_x���3�}s�}�Uf�( �,Cl~ց����ނ3:�����v�@E	g��)�x��:��VX-KNS�P4�����b�h�`���=&�&
c�ۚ�`�ܻ�R^�����9̥�9'"��*���+Z<>~R79�aT���^/�뀏~�ƨ�� ��֔�ˤ����e#V����Xc���p!�����6����iC�.7 ڿ�a	��o�1\c�W GE].��VW$�JR�6Ճ�P3��!�G3W�/�z�S�`�q�2u��;ʏ;k�F␬ys� `G��,��-#�ڷ�`�{mޝ�|Dޏ}���r��aI^?�^�Ƞ�X��f����q恵~�����6(���S�aN�Ǟ9Dra�nM/	���M��2�:c�:�@�+��U�n���B����T�����(�!����[X��Z��A�ZO��
2g�&\�f�����ݝU�l��^g�8xj-�z�x���ͳ�]�&��}j����c�M8rm�s[��RZ�i	�O�͂F�����Ԕ]z�Čc�lryFe\ޒ�E��3�;��Ɔ���R�luj�AY#4�BMJN�Eh�)�4�������4b�
nT�G�T2��`X���rZI?��d�$۩(������"���	w�q�NO�{��?���31<�r�?b̉]������,�:���I�����#�­�4�
SEF
��ݮq�KQc~Tz������(�� sB����y��ZŇ-Ӣ�f�LsԈ�U|T��bw���V�{�Wz�i�L�j���C�� 2M�X���IL�:$nGV3���Mꢴ�T���������rWR���p&N-8ۏ
��&�E�`�\%��Ɩ��'�p9m��P�e�yH��F���̜����y+�YR{=8�mSuT�n3��ͦ��?8��@�P�&s�!ҥ(����6�����}/i�j��Hp�GRx��|��>k�,'�y�y5�8�_1�F���v�NG�Q l#gg#���pZI���j�<��;D'6�"�)�T�#�ii�2nv�O4án;���6��n-�5�& H6m "��7j3b�m6����X��	�0���ޢo$�����k�n�'̧�_�˻C��e����Q�״�_6Z�V��%ϷSe�س������|+�R5)sz�3��؄_���ټ����u�g��jJw7�9|{:����)�O�r�]�?�6҈���n�r�r_E��->%�1L
p���8���W��20�P
W#x��g�ߎÐ�:���^�M��s�?��qN{�Qס�:Dv�0�7ۭ �y>�l[��4\J���R�D1�C�BR<A�-K���fa���ޤu����V�s���� s�t�����3>�	Y��ߤ�9(.G��=��y���+)9���p�	�n����}���8t��;R��a[HM�v7����pN�"u}IԬtu[��7�xeT��|�i.���/�a�^� ׊�©�zX�d��x���i�G�.��^vj��� j��RF�v���A�ݜe̅�� �H\����kDNh(cЙA��:m��ĕ �����C�I��=��t����� ��z�:��ň�M��f䜬Nu����^��טӠ�Ô2�3c�X/�a�[��\��!�{F�.����Y�>Net�ɭ�\���u�U���� ����X�J�rd�#�>�dS�a۪�%�B�QO�1X�l�:�a)?h�H�;YĻ�։��w�?�x�}�X�dr�s��0��w��#��v�N쉭l<I���妾�^��6R~��_����	���g�����s�:^+0�~���l&����޽�IϘ��^�}�q�=^ ���b��j�)��W↵�ϕ�St�L����_�:��/b���F3%we���M���C�`Qd5O^����8|vƓN.v�O�gY��H(U%>AߍmI�fˇ�<��8BCq 	��__R~9~�ɡo��n��A�}Ի[.VY,;<�rX;y�k��i�H��ź}�@�A�w�<aY��Y�H��~��G�A�S�+���>;��4�?$ttG��+~D<.f�jH�����voy��/�"���`���5�n�9=U�r�҈Q�Z��Z"B�e��6���f}�d��)� �e)xbmyޮZ��_ޏ�n^Ÿ��$@g�7�sJ�'n��1a3��q/O�7�KS��8���_W�~7��@�S�0�Π�1z�����6��>�A�P�u�&|���Ѝ�Eц!��� ��a0�P!�uoL��
��f��v䍣�y�*;�ZH�	'��d�����E�ǖ�"�SA���y��lK�~R��ߝ��un�d @/:��w-�$�����w�\���$*ﲣ��?6�f�O��Y�_8��`pF�� ���X�<��$O��Q	f�&OU�?����;��`Cht�A��Nߪ�;o�,M�-�(áw���Hdw�f�pc���(���ӹ T�H��ŉ#�_Z�������C2���!�5��g%���lqm�+�НN���9�Jy�'j�C�s~(v�'з��|&��D�gN�T�)����ȒD���ܴ���>��M0�����6{�_Zu]��P�3�9���)�WX=(�Y�[���OQ򠐛0T���-���uՂ��������r��ň�M�AgL�mpJ�wDjVb�s�4�1��X�Ud9�`ι��B��㰟��h�͑e��f־D�kWv	�%+j�D������Q�p��9�4G(�����9�-U���c�����g������6���pw�I����\���Q��������`��`ܻ<��)�����0�r��)L�{�I`,�%��_T�5u�t��C]Ӂ�i�c�:d?�it�iP�Q�;�}����T�?LP|m/Pj�*�@CY��N,*��τ�� �t��>M	���2B;�-L���@��v$C(U^3G��q:�S;R;{�	��zpv�D
U)�&t#�O��W���F :Xp�0�;�J�1d;�x�]*�|���m&��G#�M^ϖ����'.g�g��X��n�`�P7"���JUF�����1X
s���/�V��諿��T42&�'Xk!�jД� l�(�C��>���
G!L���m���i!#�Ҵ�)i��r~37n��.���=[�M�@�TP�]���v%3�l؝�v�����F�[n=1�QE.Ԯu�7��?HK����/���f��	2BX�y� V�tx&`vOQ�Dzz�d���.-)QP��}��~L:�p�K����n��_��j�����m&�J�̞&�(}5��CO6>�Oz92�|C�{I;��P��6jGH�q<���ö���}c��K��{K`�Ϧ\b��}{��qc�;7{�T|:��s�,��Դ��IK�K�p�k�kd|+�Ú�����_��x�sӕ1N�g;��Ɵ�I�T�lU���	����Vx�}��2gZ��TS=F����^�@M�51���M,�q�:�R���<�͕����ʺ�������u�o�BX�x�鵮Y	ͅY� �C3O:l_K6��׊7&�K	5]v��		�#�+�.c����sϟ?��b�hiK�o8r!�Jl�q���#�ͭBX"��o�M��a՞��Ǘ������q[���Cro����[�	2M���&k#��U�,�<�9�π�V��GJ�,��u�J�V����+<M��ξ���q�5|�r?7�&���Y�7�N���~�<�s�߼>.�����j�MAA P�1N#��u�-��,��jU��;��`�\w�(�4h�}bv&��a|� ���p�$��px�g�,��:�ٶz�!�<��}� 0�l)Q
W�p�g8�~�#&�����岼�Q��XM�Y��uYo��W���c�e��/O���Y���2v�Z�C╃���_�ʮL���y��n����{3D�Φ.�>'~�@�y���he��������Ǚ!�@� )�.�r��KD�yFi�4]��g����I;��d���O��[~ ��8#i��-��K6�0��->�j��Sg�B5���1�{���Ľ2��jkt�����J���V+n�7��~s�o�7��q�X	��m@����D��~'!��\KG�Q���eok̈́	��|�^�|=�0�{+���qq��͓[�r�8Y�����eT>Rj�z��y���y����r���hbc�{�S���Z�#�Qh�B�?��v�/�B�Ƕ瀇	��B��O���LGiC��e�q`U��ΣH��4���c��������ᎇ��(�& ��S���������dc�وM���<��"�h[�k���M�ܷp��"�Z���
��F�u5��͜^�G�Ǖ|�d���(��T4B��+�S(���HFkv��]�+����j"(��e�PN���"cbd(C����Xf�h�e�kXD����BC�F���A�c��sz��Ba�ɧv���"�[ˏ}�T0ۆk"6�H���=��y��d*��y���&�����0��7��4,�jI�/����X��hU�u,�N��aM���D�#�%9mg������;7mDl^�=վ�F�����hj;��O���!dY*�`�����̗�-:j2Ͽ�GzE�U8I��`��j/r���.���^�0RQ���a�7�[#��~�H2�R�¼��I�/Bu�O��d��@�ਬ��^�k�K�!�	��_��n0�MW0,?ٷ9N���"I�;��/4)&����LH��6�f1�a�V�O(��V����&�9H�C2����u7,t�v�Y�s*\�Z�N״��P�# hW�4��b+m�&���3`Z�Vk�е�~(��*u<�%��D�{_ݵ���;�&(i�s�]��=��:bM�̏UDUV�g�f����tU�ȥ���Z�Ov���*,Wͯ>��x\��6�Z�Y�4�YF��S��]s�34a�k��gDtŨ�$<��S^�.�,8��ڀ9�(�������e ����]v���-�D����k��.���T��t.r�tdh�d���@�v'��Ni��GT%�c���{�*F��g�U��rEm8�j!�گ���琉f�4�0�����}����>׻�#�6}���nsi��聍�D�R����.Jo>D脣/nMrn�	���*�N#�Z��C~��Z���g|(��,�V���y3��W�Ě�u.�J#�U�C�wyl�0x�P\	@��FP�ɵ�d�$?ً�s�S�%e!�=��+������~|�t�`��G�-r/J�ϩ����7�X]	�I~�BJ�M(�4�}ܟkT���f���y�qn}(����;
����z;���x�چ�=�:��m2$;1`�K �G	�y=α����)����3�o�j7�'���EZ��k<:�{����¹dg�MN�{��R��4��W��Ksa��ݤ6���=�����C��е,���l�����G\��S���w6��$8f��Ǘt�K"�O�U� �V�4S_^ɒ���X�!"���ee{%���jۯVԴ ;F=Iwd�:ݒތ�|�Y�}j�ș�rN�^��A#��u��9~᎝��:eH6���`)ݭB`�=1 �����ߟ��+H���I7��|�>j5��P3�o�I*�P5LXq?�(:��>��#�c�2�ʊT��>t6��*������$���xl�"�)��a�1��؂z��Y� V�����e)�q�#�C��W��Ģ����Aq-9�9$��B0(L'E6�{}�e����w��N�)�;j~�v5���
��'�����6k������t ڕ�
3?J �E�a��AU���~��k3I��,Ã�XK����Y�Qڪ�g���� �*qnyJ�DΧ��T~��4��� �GG���玉erH}�����#�0��ƅ�	q���y�� )���0M�*�M��IFUw|CF���|���$�9#�](�'a�2zl�xה��W�e��R�[U�᭢w��0Nd�+�-
s�Tp}/�_����o��M��.��y�5�������D��Nͦ�ܶ�s��31j3m�N?������c������x�u�-#��lӉ�K� "�SS�=���g�=��P�O_=4у��o}�ݏ���M�(�x���߈��wvY�j�@��2���È�
moA�Z�ͺ���U����'N)��9��IKgx��S�0�c��M�w9
oR��n(������}p�U+�;�R�g��xm�q���PF9��FzC&��<_>�M8���K���OH� ��w�>�0���+t��q����c�)򝽆h�������;.݃_����#�i��C���1Dڅq���(��XK�Ooh����Х��?AU�@Iħ/L�"_�����T��֘.������]����k��5���yGO��,�T�W�V����?y�Ga�Tp����C�8q_����D�뫗�=x�F��d��)�>�z9.��/�^�7�9w�B 	�����Uǟ�^߂h>,nCx8�oy�62��~��2�����X��W��t��e��oyVs����'ix�C(�6'�l���@Fj��I���#��d��� ��t���ˌ ��� ��~).E��,��}�1q�	��{�fW�T�\P�e�q�K�`�@��P���7�T�)A�Zd�����ov\f�C1�bG;������b�ٰ��3bq���nǽ'���vq���\=Ȫ��A�Ey#� ��-�#�ק�{�|#hs�P�*���2� g�X����������n�.�Fϖ�9�W>T@��m�z�t�	i.�D�c+�c\������<�.S�
��M1�Nc7y���Z��Tn��<D2�TS��k��|�׈�Q�_3�qdK�v�R�H��|�d�rȽ�Q��5�2Y�k��$|i����f9�����b����L�:ef$���f_	l����Y���/z��@y�#�Æ!�{����J�C���Q��C��2ўd��f+jy���|�:Q���*��&��F4�l��ax�tk`)��z��"y:HT�x�1GI^c 5s!�
�*����59pX$7�ۢ |�:[8���1S0��d!���ʨ��o�ɖ�G�q��e�rO`'�2d�<j�v�����v 6��r�Xm�j��ڿ����\*�u�R����ۓ�|���b*�(b���/�9���h2���\j�]�ʬ�[�ڵ*z=}�+�TٰήjDƏ�w�)����j��_]I�%q���he�h�/��@S.��d��豷<ӝ�!*���L�f�$��e0�H�HK��l1"Z�v|t��$����\�чQ��3r{B9c�2И��0r��}<�Xr�C���
�{�H\=�L�	��d��Z϶[��1����YB��7-����L����\��"]*3Y|k���C������#=N�|��/#�O��GYjkZ&Bf�O^���#�&��b+�O��!�gB��Z��־�->���793R�����9Y�^[�P�$˵��i�����.vHPW��Fق��_4��C�"�/=j�|��m���Ԃ���7K���eNdH��$�Rh�D��d�[Jj�a���=>jթ�Q6�Ĝ�{�{�[&��O�}C����V+43�����ۃF�`S
G��!����5�N�PS�v2�#��@|�=�^U���̙�G��bn�	CE����:���*g{�� $�O�d1��֌}d�K( d�2�G�ٲc�Q.��<�7�>���� N	F�uI[!��xq��N��6�,���έ�2;��80kU����o<��"�&�7��)�4�;�U��/�6�%̥�i2r��i�V)>�� S*��ǭ�O���qPZ�;��,����ϼ ��3�%4���VIMvͣtbb��j!]�z��7(*|�M�=�������٣A:����A��6#�j�a���P7X.+�����}m���[o{��RG�}���`|�>^�ǯ�:���Fw���
�j�#h�6z�9�td��`����N�����ŊzY�q�ȷ,#��f���a�/�Er|4�5F��dm$��%�
��;.P���V!!�J!�MF<��M`%-�J�ٷ����m���-��a�M�g8]�ei����xC�S5`�}���{@�Q4
\�d!��jX�&�^���Cؗ�j��6(v(�Y�R����K���x<t�A�����z5i��c	���Wt�[���@� ������3!����z���7�W6^�pKXA���˝�-<�
�
�̐��>�� ����'��0s�tN��F.�1r�!�lweQC:���]�'@G��IX7�
_Xbo������- 2l��L�c�~<���7%�ȣ�uA�������	��Y^����B����YV�-=�Y$���N�ey��^0�|Jt�0��#TZѮ��G�a��-�����r���c赘��qi�Ɉ	%�o�r���[�x ��E���$�_�,�'�&�f܀�lA"�%Iv*CWDϞ�L[pq
�Z{�֯Cm�7�p8I:���DK㚂���ǆ�*��{z+Q�,#��[\�\p��s��j]�[�$+�&����
58�t�Q�gI��4�E}A=Ō�f��s�G�?5Hjb�mCW�ٗ�sF��T~O�US�8���GJ�����1kSMη{��ΡۿiA+?d��k5���[�Qƣ�k]��A��&�%�B�j�kP !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`accnefgpij�lmnopqrstuvwyyz{$}~������������������������Й���]��s�����������������������轾����è�2=�x�
d�>q[5
��v�S���űH�w��d���*w=|�Ȯ^&��|!Umy�;���l��]���<�JO���}r��i~�sp�G���w�H�J��\���"�H��|�iz�-��}��z�ci�.q�a�H(�~&��q�z�V�g(%��c ��M�]Q���ݧ��^ ��5H7��l4)���_����0��z��	��G�,Y��38."@���a���M@c�sy����]"!��
e��q�=�a�KB�);H��"��X�:�x�����������rV�5��|!�ЬL�Hw�"�3vq?�2�n+Ԛ���S~q��}��%����Hɍ
g��:Q�J�թ��>��9�sŉUzANj���O���O����wI�DT(��0��U�@� �X�0�a�>�l)��r2ӽ"~j�n�t3�������|�I� `��ӕ�`:�qE	�85}�d������L}Q���0!��BЌ�`�v� �\ҥ@Lsݼ���{'���z���r��AX�75͌�H�Ia2&��������	�wI�����s�`�E��c�����;�#0�sgS��o���b�]���:�����E���+��m����J����!Q�\mº������Jc}U�z���y��n.'y�<��t)F*�'��d��"�n?N-��R�IB��'�
,���^jA^��*>%P��CI�!�-�z[=�d�)�w*��� v��C��=��.30�s�Y� �̈́��{�狌�X�x��8�~��Y ��/���R�CO��ĝ���aR��d/��%�[���g_j�7WV�iZ=��1��9�����lY���\���v�~ǋ�M �e:�/l��ˮ
��C�d�����)��I"Iu�_!q(�&���"��N�v�w�\L:P��ٱ�!�o�j)9*�����1�{r�y��
q�CK�yϲte��e7���gF�ߝ��6�	6�kk��o\ >2��`r@�ʅ�~>S�\g�,�F��W��Wdt�x��J�*�kM�L�X��-$��E�}b�o
1'��磭ǁo/��먿��Pۨ�DX� �bC� h�I}����ub]h6n"��`64���j��>(�Ƀ�D:�s1ts�CU@�ff��QIgJHMb� T��Z)S��Y��y�ΰ��K�TZc�"lCB�I_p�8!^��x��!��au`{'����ԋ���h�n`H�G���Y��������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRS|�VWXYZ[\]^_0�bcL�fghijklmnopqrstuvwxyz{!�~�Q��U��Y��&]��PA��GE��}I��oM�����������ř����ð��������������˥��PǗ��������������ԔԐ��������������殅��������������������k�WskwaFii{ffnCxzeeEWP{mjr]uq{]UGDFVV&'(nO_oBCBQ_V][Sv89:~DTJo2.!&76FGH/?9/=$$":39XYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~�������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSVW������ހ�������㰥m�����������e��#%'%#m/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomc�gecs`�me�l�L�l/�F14,}SWHBQLB@DIKLI_FUPMFCahv�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#}j-#i& #�k%'%#-/-#�''���������C�������������������������#%%%#)/-#%'%#9?=#%'%#-?,#%#%#5�\cdgecmo}cewec}mcewecmomcugec]_]#%'%#",#'%#=�=#�%%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]o]cmfecmomcegec}}cegecmomcegecs+8[Q'%#�3-#%7%#=!=#%#%#-/-#%'%#�������Ý������C������������������#%'%#-/-#e'%c[\WD'%#��-#%g%#]�]ceWecmomcegec}}c%ge�Cgec�]]#%�%#-+-#%�%#=?=#%'%#-/-#e'%c󭸏����������������-�������������#e'%c-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������Q�ʻ`�\��0w�R��vU.�߁d�1��U��i0�X���LY��k���hXБ�D?qf�#�4MO��.�v���co8�h�AO��c,T�JΣB`8�=j�G��������* �?o���P�N�Q[zs���(:���/����GD��\�01��!�E-�����sah�&�֑1dQ0?,��.���D6f2y+�_��a\u��� �w���O��_@y��Y�<6?TTѹ�"#ꥑ�	`7_�E����+UoxH+�w57�Bd'��Q�#�J��ws��KR�3�}�y��e�F�e������к��i����� ���p]L �J%�ǯQ��Io�_�(Cͥ�Ȋ�/9�y���9�>b�Z�I8�!:[[Oa��*|'�|{����]�Zݠ/��:c06Z��P��"JGs]���1���������h��
B���}G��9��~�_�6 ! \���7h�4��s�ژK�1뗅�rQ�����ކo��#7eeiHs��:��d�!i/��)��-$�	��!�f��!�˹���!V{ќ����䳘1#-�&�!�+���v�i]Pr�\L�	��.�jm��7����ؕ�Ei^	ٚ_������l��������	���yO�.�Q��dV�=ӶouR��?٪}SBfR��s1���_�Ŋ���Y^)�O��7�r������P �v������i���.cW~��Ա^�[�k����6�op8� g�	�ѡ�������B	*���7��U�m���pː�.�%�Y\�U��l���_q���bV	� �\�ͱ����Ś�.�A�Oŏ �~?�4���\�*�0�Z|�mD*CFH���Ϸ, ����
t_5 �K5��J��z =W��T�J��ՙ �\��t��Y����Q,�^F/̪F���;�N�� ц�c�g n��!q�.�H���$1������|��K���o���.��[����h�AI���<�7P���A޷�I{���|{�PV�׫�Yf֦���zw��6�I�ZI�PK9��\������˞%����(⅀Pe�����,[����TÄ��4�{�*:/���nߪ�OSv�3x��d�4W����i�M��T����qR˜�U jc���o!o8�B�Br����l����6��jϴ�ʨo��k�y�G�X���Q>Q�vpg}k\�W#��S|s1U�y��iܸ.�Q)�}�ݩ C�'|�c'A�oa��]���˕�j�������d���MIì� <�=*��:��"���6�i�s�	C0��W=ɽ�<�P0�g��Z��%��)9���,�?fz�i?�짦�(`$s������|�N�0'a��� �ke�i�v5�i6�-�%�R�@	�]`�KĻ����تΫI�s���|\+�[�ɋ�L�\��Ő�����Q�[_Q��1?ʞ��h�]�%k�P�fA��g�3���,n����vBX�v����
3H��f�s��I������m��	�x�2��(��ז؟���U%�捹�V��� ��J!��'��?01�_���d��?�fS� 9�]���}Q�[1���z3�59�������I����A��Wq�D"�5�S�|���>�m�xT'E5b�	��N����j/#�g"����a���c�U�z�Kq:�@��8�;6ԫ@�.8�ΐ�$Wz�����
��v��NJ�-�"����1<�Қ)��������"�?-���LO���L��
�B�ħ`'� �U9�<�}I��У�>tж2q1�@U�����y4�9�Mi���S9��Uj��u$S)�_�蝻W�I�s�<�������R��|���9�3x�H��^�Wᷡ�~w���c4���*E������I�� 5�]~����g�
0�#z��TI��F($���U8>b��rS795��|	��V�6))V�3�����+H"46β7�9�vP�0Q���k��v|=¹��VQ����
��˄k��|ڀ����P�T��Sz��F���1>���r�������� d���W\f̋BO��)����kp�����z��NijJ ,���������e���r2Q@��>CԺ�TO0%�ݬ4�<g�P���%1;�N��.�ڝ�K�s�.��N�z骡�s$+q�B}��k>H��VB���I�ad{\H3����t�C���k�vz�$),�4��v�^�{�z��>���������A:�*���]���]mP�ݘ��7%��� �3��im�B�+>���)�#��r
����}��W��i#B�6����F�H?iXKPe�<֧���@��:�S��ȫK/�.%��d�@P ���6����λ���zX���bҭ*��$tE��l�y�U�	��h9Ӡ�_!���\e�&(�x>K\c�%F�E*�c��~�Z�Sn�y�(�<������>V�0�VW�љ�#�m��X�
3���!ٮ�j4��3��
'L7j(ނQ���u.#ً*t	�6/6����0���2����ќ.��ʞ�&���7�xo�J��D��|����r�Xq�����=��(��-P5@		y�����Bg���D�b��#�V�m�����٪�Ve��{��V��Ϣ��>R��+�B�3H@T��i]m�>1L��}���ۑ�e���=�Dzg�pJ��T�SX�-9b���iٹ�Z���͵�H�Z"�L��(����)���!��!��D�x�MУ�/�UT�@v���\,yа?�{���%�ՆЖ�%���;�t�΅y
��yh�֌G����<�Ss�y��U�,���ٷ^�d��?\b��ීC�Wi+���:k���?v����A&������6=�G��6�,�L�Co�\U!��$?�j�/V\�s]57�Tu�u��F�3�-m��h���H!�S��������F�ׄ�p�ٕ~q��Ucl; ^o�� A9�@׏\ə�|y�K���)
���|�s��������#�h?2sg����)�0�g�*���
���Ff�SU|�_� �$O6��j�{���S4d@�{�㩳Bd�h�Cyy�>�/\Q�^q3}~�2n���>|СK�-�!E[qf�u�&�	�0��6;p1�;�za�����v�J��%r�y�YR.����V��v��Q��3R������l�9���� &#xM�%����,+@��O,��1m�q��뎷�21!o=D ��-X�vK����L�Gw�L���sm�Qh.��cEN' ,+Ë缵w�7x9t���s����+b�V$���,ꕺ��6N�� ��Z�̠-�� �ǩsZ�.F�KR��0��lU2�LP����0����S����.��	��C錭0�q���:��U��@�J4X���jy��
^����9+���

�4��E�{[\�*/�.$V4�@�)��{>,m^�P4�*=��SGM)��9���*펔��I϶�+y='X���)V%,n��jT_�Y�r)�R�JRK�="��:�K��(Tª+nC�˗�ݸ�fZo]tT��.�T�;�`h����G�7qL�*�o5e��	�jO
�dy��n�	������I����U�S�9H.��6��2u�M�t��~�� �y���������'� p�-��a���U�J��H�# ��l7�؞�����#�9�.�:�muX,z��D�J�3,h&��c%գ��;�m%����\Z�1��UunN-U2��s��'�!7�Xǃ���?�$W\r�(����2$S]s���B���a�4�XԚ�U�	�/3���) C�����WO�0�5.4���^��プ2�@mC\���lWHu�_��},:����e�k3�.��/���ue˭1�C�+�'���"w�+�ߗ���P�5���!�����BZ �G���a�$$�U��c���v[�i^��~�9�HLrZj����s���
g���/Hѥ��ȿF�~]��E�]?���+Ɲ���W�P I+����Q[�`�tf� ��8���|�~)2�4C$3|uҤ39��W>����٪�m&v����M�qv)W{����1��\�C��K����}G��2���{/�Yb�@����յʻP��3��~�e��,��M��)x���,ղȱ*!�l�\�*�l(_\��� �]M�Lz��3G���iL�#�0� �p(���-B�J`�a��q�g��ٔ��"_�!L2������DG�'����}i^Ăj�S���(P�D�SzOTjJ�g�n��+��4�8�0WdC�}D�S��,`�%���)f!R��]M��-%���8�x�2����닙W̞8ʣ'%#��/#%'�e�]ce��Ē;`T7}���a�����/ege�h�.�'s�͕'%'%"��*�R��+/-#D��'���#$�1�.9�h���=R�q�'n���������^�!�H.,/�v��*��� X/*���'%��U���fze� ����ﵽ�	������A�dN���=v���qSw(��bmG[w�	�!�5Z�-�̖���pe0��m�Ҁ�d���
�0������a�$��Tf���)���i��8�\/R�F��_�%Z�4WǄp�o�rv����"c!G�7�)_n�G��**�Z}\���Gk~i�����Hw���n�}~���+�3�Ud���,��լ���N�z�8�O����-0�=<ҩ*/lݞ�>B'7!]�4���!�wB���pK��oXt��BW��JLq�#6D�~?��f���	�~�L?��T��4�����������b������&���ϭF�V�����7����n
_�)n�0��Z�JI��;L%
�6@%���<����(5�R��Ւ������	<��8
��A�X���Y�XP?���Ή.���x��WA��s��cF>�"��O#�������T#�>�x^ބ���1?{P���}�������F��%��������Y{t�Yv�(s�k[��Fս��Nʠ��PW62�G��T�Z��d�,i�}c{Z i���S��B!n��}�4�9Q�-��γ��Xc�R� �ֵFޭ� ��S�Ai��L|]��&�ڙQ�Ф�s�"'�=;#��1 �"�EnI������9&Al���IP]kW��; ���'�jj$��cj>b�8K�X��,�����s3�Z�6X��^�>��]z:0Q ӑJ8A�B^My���[�ѺTm��q�hl�k$�H/GϽ9)k^���#�<d��
3\��(�V�-־dyʎ��/]���l#V��;5C�C�QԲ!G�j����`�h�-N>�+�{L������_���;� $�Q�>�������  ���ޣg%\­oO������e������	]�f���!�0�x����f���)�94��֞?A�#j/DG~:!�Z���< z��}ބ�}c?5.����w:i5��<��	�rܢ F/ʔ����YX�#K M�*�Yf�� nu�v�	^�YO�E�'���C��~j�f*��8�v85Z=+���5["b�W
#�BR�����Ѐ(���QR�U��ֲ�Ƒ��_�̩��	`�f�:{}qM��4��tl���P�E���F�L�&!�z)�>"l�9Fr���)� 2��@��iU-Ft&	g�HSw���A�6�bAk�?=w�&�­��Vy�O=�@�"S��ruiks�Et�h@�����ۄ�˞<�13������ǻ8���]�^��Fi�Ƹo�dOjռ.d	ECLN��N����-{�u[�*�'�%�� e�3umИz�~��e����,��q�mr�gF��9�&E����4����s�`���iT����/r��>ߦ�mN��pjq�ˁԀ�i�]�p��=P�Zw�v��r�b$ӅQy�#�`qaS̙@_�ދ�{�]���`d��i�K�X��
�f6)�0�W�S.!%������58����k}~�1J��1��t.#UB30IN��?=�`莉�)�����T��P��az�?�('���9y�<GP�W��"U�H:��]އ?�v�n�Yl��3E��\�v�ȃ]G�9(F� j
��eg�>��vnM93�d��٘�*9�S�K�Z+p���$c�-�g��b�9(&MBXgh��'�=lѡ��E�S�T����x�俛�D�\	$�2�q�&�am"�`+{.J���ȖxK��2w��B�Zs,�����۴E����2�M��٤A�8�k��{���W/Y0���y'��O��``�US� �2f�f�K�H6���	��}��ގ����ZX'R?��}���:�;Y���^6�Ĥ��M���a�m{����O�D�����s�hb�1H��o�L3<� ~��A��\M>Q�k����$�*j���몲�r�o��ʧ���_>��� NT�9G�}�І��0��އ�a�o��7��_�4�V�Gc�����?T�6!��`�z���/�4��>�|�!��>f�5��:hE�ݵ���<YFM����U��bN���ȁ��8�OA���9M^EY�By_�\}�@'z�r���A¦S���;8�&���(�C6��
�g>5���Z!��>z�]�T��� �C��c�n��H#��Yy@�6̲�*��4f�ԑ~�}9�+�c^D�I�c%�?���f�C�7c��n���*�ql]R%��ɯE�w�KcSf� 8��(KM�9����K�E���_Ft��~�g���Y�N1�Z����T�;�C���l�-�.J��\Eb�nZ�f�6.��T�Q�9?
�ٿ0�ny���I��D. !ٴ+��K
s�Z���i&�W�0U9k[þَ$��Fa�hOwn�z���d�צ��=��;'�@N�i��xz�f��Mb0����G~
w�!@�7�=}���cm�
.&`�/I�uzW�Y��H+�l��8���.�Dq*kk���U�:����d0=鐼Kt�[B�e��Af���n�^�xl}�����T�#.��5CW[�����Ӟ�<r�#�!���(l�-"�:�iq@ޭe��Z��u��a=Ɛ�W<��eg?a��7��W��𻻚��?�#�9?���ͪ�Fc�>�?���S�9�a�����y%G{���4���n����r�,6)NA�]��;��aH����)�W^��m9�:��|�D�,e$���C�c�禤,/I��c �z3���p���H3C~�`l���|8���w�`��Ok�3W���͕��/�wMG��:Jc��C e�]�($+���C^�+jOe��4d�ٸܲ[Fq͈��ے�c���N-���s���(ا��M؟�1��~�cW�&F������p��A}"}�ÁNZ�gβ����i�	Y��B8f��v����c��1d���t-�ى�(k�	�C�.k�ٚg�Ⱥ0�T�o�Sͽ�
�H-�����>M��3UL�T�-҂��=�(;U+��jϴ&�M�p���8�����,o#GW����Sv�Mj��)��+��;���{(UR��Q�9�e�0��������
�R=↉�^#v������}���ݱ��&޳<݃�~8z�U$��%�[na���H�G\,��Zs���/����	��]E���H8H�љ3`o�,���4!��ұ�w�X�'�>Z�WSE�o�j���Q�ܛ�{0���c�NY"��a}zJΏ�T�6��V���'T�@���m��nJk�W��eH��п@=
���F_�%;�\&�LB��Η� ?�$2R*�mVzUu3��H��I*�☺şM5v��
���Y��~7<Pݹ�׵��AQ�Y�T;�җ)���_oh��w5ȶN�U�AM�b�E�$��B<L�(���!p�Ԡ�i�����������*��d�-�{ˌ����B�_����A�g����ٮ�1a9)��>^�IW(��Ĥ�����zY��=H^�8��up��A�\B9��"h��LEp�����J�D.w�i;�w�v��K|��vG����؅�r������$zܠ�M^�*#��(I���z��d���3��IT� _�/G)�n/6�:�-"/��e�䞜	� 4��Y���6֒��;X(�W0ǑY��ES�k�\L�s�El4��p'r����DQ�.MIY�"3���(�j�i!�n�?�#�p��(����#h������ڬ�`�`0��d?B����RJ%�J��}c���f�O���1=I����`ۿͷ�������l����` kM���@�����⧥os����>]-X~��-�A�*�� ���g�������(��BĨx+���w�S�����1�pm����A_T��JVn� l{H+d]t��� N@$c_��;��ηA�6�K��r�)�S��>�p-��f4��ܕw;�et*7�na���D�/�d�����/P4E��9��O�o���JR���^L�����w��Z�}��c$u����VkƮ)�^�T���Â���ƕ����0�?h��!W�H�,'(@�$��P�%�e�wK�"�4[Q!�ƱV�x���r=k
���.�lȢ{0yK�^�b����
�v�4Y��sj�3��A����� [�$�6�y�ӛ��B}y��\�+����)�W��*<+L1�OGoI��o�̦xs&F�w�l��7��/�1��J��$6)ި�o�4� 4����o5G�M
�;���C~M�O3V9���3+�W�%sj��?	3���=:Q�L ����</y��%C����7����D�db�%�(I1���R��[��},Л=Yę ���	�� o1'�Z:�zJ��%���Ž�p��Vn�A,r�t٬6��Fz�o�a/��Z�j�weD,���x����e���`��ɘ�Bǅu����M?)i�o��҉M�jF�Z���&�������OW��������������Z�j�뤛Iهˁ�4������݌�[�8{qSΌ4�j>�3>Iu����^�{f��� �,n�0�a�X�k�X�z�U�=�][�
���s��O׭����H�+�6���4����ܟÝ�qD���عؔ`��}f�f9��ԛ*80@����	킡/��B>���Z���*5�E�,E�"�.���Ug�~cl����	�`�(l�"@1���|�����I�����I�e�C���	�8��j]{_vT���7n�*ף�p��x�>�u�@FE�ֹ9�1U�O$Q�WBoM�e�*0;�Y	e�#r�{��r	����u��q*����j��UO��G������ȝ:t���;����L�]X6h7���D��j�a$��|A鑐8��<& �0!U�4ے�L�����ը�׿`���V=K�(���.2?X����>�'� ����q�ǽ;��M�9�q��AzI��30zW���|�t!k�^��(=�Ay?��e�1���a֊���#4H��G������HQ��P ^�O�#F���^�&e�9 GE呗ㇲA���>Uǳ�3��*��`y:\���k��}�"��|�"�J��#�x񓌺�%�EY7L����Qz�t�?�y�ƕ��5�"��Xx#�:a\���ϰ4_��B� Í������xҮұ��;ܛ#,��,`I��Z��
��+EϨ@��/��Dmm��t�����	>ă���r/�i�q� ���(\?)�͵{�Aԛ<\D���&6-$�u�&lqq�
(����bl�W?[�W��T0������&�\{b� -: _+\==����k����2:�D���۽p�ȟA$����+�@��,��u��!<(7
����2jے����N^4�R;��F{V���dP[�����'�c�G
����X�3�i��`��DnN���P����0,ot�����C�����=�X���_tE͊-9P��N��Q-`�Kl;_��S�BN2\ӣ��RqKkX5[XJw י�:�ix��I�Ñ���^.K�������������7���5`/bZ�|3Qʫ_5c�J�6?��'��W��~ �[u�@���?K��a`WX�����hƓ�2�����L~^��S���j����D���"~�H��*t�
q�TR�x%<�����u#��>%G]���IHr�8i]e��%*���@�މ)�'�Vξ;����W��Y�	����C�c��J@�#,�Q�)RT���~��|��RZ��']�Q�<{ϳ�J[�� lE�����9!�/x������z��Ԡ���%��U̓��[�V�C����/`j�!�����G�Mg7��Ӕ���/�t��m#�����s��'�<�ױ6�̾p�j���,��)��ٙ���s���P�d��R��+&�g���No��%�%��E�P��� RHθh�������=RoR{CQ/X���R�~%�ZwG����D��f�M�$��ւW��}u���U����k^^�W6����(��)��%c[,{���y�*��$>����{f}�>���i�-)Y�J���4'\����2�&�.	dҼ����g� ZF�ɮQ6m��S5��f��"E}�׀x���>Ɏ��@����)T쀳�� ��p�'������D(�V���bD��5�X�`���	w�276B�N��R� �f�}��!�Т�QĂ������ɻE9BõAH�>�P����w4�]��L�>�xȁ��+�LP�N8�N�����,q���-�ɼ��z�Q!�z�W[yR����s`҇���QU"���i
8�p2�qn]��;q��$�H��h��� +R?�3��&9�T�����_$�{=�����d��+���2���(�{ݔݣ����*i��ޛ���r��$�w$����ɸ�hq���n�T��N���z�Hy{.���
��_�\���6�ҷ�)��lh�YMyܤ�p"�}>��]'N��&m�.�����{	7�ǐ�H�g{�[?�v;ȗ�(��Z5~W$�B+��~F ���iV5�*��:�gчR��^�"��d�\ή\$�q���mlțB�x��Z�|p����\uv)����H��d,6��$~�Ak�q�@n��T��=�,�&W$���},�4lx��Z����@�n7P_B�n��[���C"�6����!��r$����v�7��� �,�M���M7�mu��Dy���H��H���s�W�(?e���hF3+���z�{>���&}�xj�_�h=5�|��<0Q�QX]>d{<��Z�X`<	mǂ�i�R�k���7�ڝs��+Џ����-k��j�aB�DP�'%#lB�8e��f^�����=�$�W��$hqP�C<��z�4wi��������Ŭ +��nou�����D�5�^~9 s;��}47`�7�9qHy!/���b�`P��|���Px�^ ��L-���!�S����H����ihVW[���i�~X�j���r��^�c�@����`�wE�����Q�:��S���to���TD�x{{��zҝ�M��.�Eg�^���g�L�[q�3`q�9:J�Lg/h���N��̲-�rg�}��<�m�Ȧ/#8�Jr
��0��
(U�2�@=�*�}<j.����FZdm��Z�ٞ�ƚ<��:,�z�R��y���M�M�!��WP�=k�2lAcqO�>���Hg��;`{-���l���p��\�|�au�8&~�>�oVs\M�-bh1W�;�y�j�����K�4�����ڪb璹�tJXA��0�^�)I	èZ���"Ǔ(X���C��&��Clҥ�6�t�����'F]"����z
l�5�}@$).P���8%UIQ0��(�6�u"�R��L��@p�V���]�ٜf#<����T��N��G��$M^!����#S����+?83���T�WΉ3RB�(�X�NO��.&e��{s��^�pVf$A+*x]5-���s����J�J)0�O��W{�s�� (�y1�! F
������99/��C�w���TDHxc��?��#���5#�M���R#!C2J�Y��,��B�mw�[���%�x���#^ϝaŔ�&�fy�PO�vP2��Ƣƛ[������NG��T���D��E"�qΖPo3��^�&j�P�����4�tf?�9������ls�(��1j�ނ\���_N[G�}�xJ"��/U�c�D���nY��p��˻�����ڧ�l��M׀Z��y4�>�M�S#�k���6�;�Z���d��ϽI�qAvqʬUލէa<��
�g��b��� ���-��X�r{ɢ~�8�#�-1��n��`�x
���T_[��'�Yz��늷������ ޱcr'6�A�E���ۗQ׀V�C\Ni����� �C3@&"Z�;a�l�����'�ᐵ�<T2u,B�6���*.�j�wfox�*}���r�>}��5�����b嬓yR��YH�_�N��r�	����;΁ ���:���e=f:�Є*���u��Pݔ��|����cvȏH��3� a�;}��s���J)�ҧ.����Zxѩ\�1qx��@��t��]P咺I�#��Z/����6�*��9$�6pۃc>�;��ji#����)M?�#�����Y4��.w�[��d�ݯg�_`Y����� ��4��u��S��M(�ُ;lR�oIm�W|�� �6��芺*v�uF:��Ȱ���~|�]��c궓�vӐ�bݎd�$b�U�R[�v�T����YNx������(�N}:�����ig��mb�<Ł���yba��KҞފ܆�َ����m�U����/��I0�hL}%����.k�?g\���M��|�yD� |Vxm<iv,!;o*@�	����~�aTW��+�]ƕ�ύg�%'��]��=K��Z܃Ly��y�r�ʪP��A�"L�-�@��5�f�/���� WR���V�2z���z��Эŭ��L��R��i4s� ��>1�~��7���W��ֆ�c�W�-� DvrGR��ɰ����.;A��Wt0k��Y��8Q�Q��&a<R<E['׾������p��أ� ����/��}���{�r�O�&��l�)�KKj9�`�<��!SO<o�z�4�5Π�1J�keT���*���-}|�BM�<'�p���Ӿyx�+��3g=�����d�	�ԑ�Lzѝ��Gq��D�BF]��p/��}�c��}�]���ˢ�`�X���򦇔$��EW���m� �Tl���n׼�t��r6$<L��ު�ɜ���7yG�:ȳa��$FR����)IBgs���Ol�^�}�6U[*gĭD��51�2[�	u�sܗ�6"D�$x-�l�뼗݊ҊI���	�D�8®ɮ,��	�u�E�(��ժ���"׸
'-�#���`��_�Y|9g��(1���P���S���4E#~Z��+өN�%Q�N}�4]���x���P�Dj����t�ِ�2mT i�ͅ�@�lc�>�ٓ*�Xsb��4c!��8��9cF�N)��%�����gӦ��� �hl����dM�����5*f�R�G,o����^�<���N�rIf&�����$��y�X�_�ޅ�%�Dz�ؤ:�U��$.5}�YK#I�*��'&�MU*}�MN|l�ǜ�ܟ������}�
���Cp'�Kۦ�#�E���7.V.${��뗖���C4>�Ɣ���Ŵ$T���CM8���#��F�I�$�v���O��Qu���¼��?��6>�?7c+�D�SGi�ȓ;���I徶��Z�V�_�z��~��@��Ok׃�����,H��"o��s@Rå�[U��K$!���٧ag4�馧m�E��粷Kkj� ���!��*�(NFu��6��
Q(���1����qs`��͓�K�N�i�����VZ�6q;�gs���Pc���+�L��ك�J�q�m;�"	�K��pN�����볨2����'�M�na�<���R)�8c�e�{�d���9�mys�3ȟq>�B�\E��dE3u!P:��j�%D�81/�p!�8A���d����3��Ч/� �Ռ�x2H�����=�lY�����v���侦��U��uo�`��Dz�i�����A���1ȹ`���4}(cù��e��udk��IK�3�E��qbSl4�{ �q%�7�s�����4+޿5��-.*06̋��}nnb:�j	�<��b���8��vKU�XS�t�p+�9��3�ۤ"@���h�����E,y�:_	�[ِ���zi3Ɋ6?�@�Z��g�yx1V���<�x�ip���*��tS��z��B����8(wD�h�V4����N�#�"6:-�QD������Q�P	���U`���/�)��^�3�Y�=�,��,���M_�'d�G�[����5���!����i�+,P��rȉ�E@�I��nR�1y�d�R9�/��AP��Q���%�g��\����C���N ~F�jʏ�ZGKr�iQu/�s:�>�D�&���dU��g���`Z7�XDZ�k����<?���-�����U�dL�I�%
��H��r�Q|��2���}��vV�K֒B��9�D���^1K�VW�j�Y�ʆ�� -M�%��v�����]8�6=1V��}�=�:d%�Mg;���,�{�BOz����$�;�8a���H��۪*Б W�ĵqt����xG�0�B+�D��*�t ?F=����ہ�=j\���3y�씦݃�aa���/n�i��(<ȥ�e��r�;pE �ɓ�T�s�����` ���[�,��prRo)A	�L�#��j�~��W�sl���_ԴV(��#;}�~'}���V$����Q�ד!m[(|Z��٦W���
�rr�:[�V�lɈp1=��WW�d��	��a�f����32/`��8����>�r�� ! ,�v�y��)0�-���lE���9�pT�엲��*}	B�,��ϵ�p�γt�8�� t3�?O���Qqf�0�˽�;S0�����ܻ�$4��tv�Avw�'��K��y]g9.���\᫖.��/Q���w������6��p[�=�;.HԔJ�2O��2R�e�j6�R�w�/��Ζ���� Xd�d5��[�����F",`�&��˭�x� N�_�v���2g�'�J�����q�CʿDR&x'���J�=ߔ���j��Ĭ���F�CJH/��u`�o�Q���mT��-������ɽ7��*ө��%�QL�%���y�j��)HUBt� �G4�/0abvL����&�t�����23ZL�(*���U�<�-e��^Ib��o��q�
�giz4���5�;��14�)�Lʑ-}��\>�D1��\��r��e:���?�>vw�P���9�"%W������=x����G6��U}�;䯉/�vݢ�����O]����������Q����9�o�l}�`Ϟ�Dا�&Ds�y`Bt8*�14�XJ3��@ �0>�w�G~��jG�Sކ� A��_os�B�M�UmkWa�4ŷ���#�Il�GP��r�j�P�"A�+.۝��1�~  FR��J��G��2?=�(��be���~�7�fn��,�Y�1�j |���(�;���=`v�,�� ��M�R]���O�T:T^�!�((1/e
& ;�{f���o����. tR'�Қ춏Q���pJ���}$�i��>�-�C�v�f��u|a�s��ߛJ�8�w�b�o!�I�i�p ���{+ٲ��.2Y�iin���x�i�&W!��u.��(;)�����͹.�|{���'�������L?�֋ɑE�`솬|i̙4@��^��Y�T�)L�s��NX]���C���[�r�����A��`E ���li�\C0��WI�օ�\����u\B���Ug�9oy��[97�;�i�WT:ƣ�ԏ��Х�n_c��3������#9�La4� j��˷7b��VBK��x��H/P�$�mMϫ��.�S�[������)��;G�e��Z�����K����oR��6����<��G�������Sy!m�_s�S� n�a��9�����E���2�3�e�X�)�4��Ę��4zsu�{�@0���$���g���Ğ	((0>ᗲ�Ӡ�1j�G���V�ō�L�u?��6�Va\��2���-V
!�lf�c�	wM�#�^d����~ڧ��?��\���aKE��%
�b�ܧrŚOf�	B��Ұ�H��:��� �,�6L�FY!B�_����
	k�np�{��e��(�O�F�*L(�C'x�{#ͪ��y�=�
��Qƙ�����2u����L�h�v�_^�Q��7�Vs/Yy��\b��ӰxB$�6&�n�'[Ad�b˂b�%s"|����J��+�cT��B�ϳ{hy�ﱌ �ݻ	6!r�2M,ܢ2��/
��`ͦH�)�χ��Kxo�] �F��e��"v��=�]Znx��C��CZ3��_�_X,��Oq�H��mRCl\���R��c��*_,�c �S�%>��o�
���4N#`Z�1�y{��H�t���p���p���I���G0���h��rfž2��(�Rp��Af�HiR#�=2�jGWh;s��$$���h"W���8��/�jjO/	,�s��]2��lۗ]L�}�i���L]����Gh��	IA��R�sS~tf1"]�����6P'r�7��{c�(�y?`����`�������1i^-���&�����߂R|�s���0!��{�ϥv�(E� 50ϙ�����1vAie3kg,@c��*�(��9\���{����s�����WrW G�'�W5��{�0Hu_���rw۶����K�d��Q�lNE!4���"���;���s&Q6� �-��J�����l<E�[N��ӎ%�]���q<�����^�Fu���kk��?F�<��Qm␔»S���79���|7}�����>-�G${ٽ������		9)^�����H�� ꥈ��s�QT��Q��>���8XpDԝ��[Fl�G,9��9P�	��C\���7w^.�݋0�/M�]���3�$	��������f�W�La���s�2�<L0�>'�t,p*��DZg2/��_#&�L�� �+0G�V�n�R`D�#�{��(�*�u�mXN'.�a\���(eg�u��AX#�Z'7ghϠ��a)�!�c i�J���,��Y8j`t*_���S�4�B#��O ����?���f�3��4�:E��eZAriiHʠ�Ȑ	�*�M�+�U�JW��3_yCW�~��Ƣ��';ws���YGF4�AP�����ɺ�-y�߶�Ҩ��}�<�[��
����`��ʸk����_���Y�}d���g���(�ySQI9dMY�Z��S/��G����8+�`_��| �����7z���Юo�8�i8�]���C>�^�±���"�A�����I+����j�%��E���9r^]��t^U�C��J e��z�2�@�j5D'�2���ڟ�3O��H����<v'�^���>�?�@�c����f+�E\9���:s�|�I4c�*49��j*�_	�M:&���`�~Wb�5�&䱚�H�ȶܿ��;p6�׹*N��5Ϸ3*)�I֐l<�8bJ�kh�=H�����#�\�s��+�L&b�5w6��g5/䢛���Q��#�aB�QD^x؁
�k�b��L��s�09h�$�
��ELx�s���*���3>q)�;�N �O��0���#�_�]h"�o��N[G"#�TbS|<����%@������4�c�T2+�D�Pފi����LTb���?�a��R�.�s�u-KI+�p8�䶩��4z���^����4�\��\���� A�}�������0癯�Ue�15�o��_�#'6)����z���JU:A&��[�k�:`�<R[�  =�'������sk}"���}�1����]�R^\�"ȉI�E'��Cz}���ꅰ�l��΍�����}�>���,�%��L��:F�$X3X��ي����,A��5��F�ұD���h�a�:�WT�����NP���6 >�__=��B2�`�<���*�ȭ�9�Py�%��D��z�R6U����,��!�T$� ���s\M��;(G{�0ۛF�HO"Xig�GW��2��5Ak�j6���'KrJ��������!۾��n�T��f6�ϙ��N�MX�-����� y���D�s��L�j����xjd��J��(N"��S*kW/~72H�LU�1��4���V#_�'\��λ�r��Δ?͛�G�H� �tVC*�4���$�� 6T}b�f��7l¬�Wa���cA(�&*ơ�l��:?����'I���A�FI*��x�3��W����6UF��܇2���;������8;{`�����y�z�Xԅ�e�Uiy.]���'�xc�m�!��/�o�Ho�p�P\wY�f��*��HW����hL�ߌih�@BX8�ů�	 {9KƩ�9F�ό�O�O��Cx��Z7#I��D�Ц!��Hi���n��b؃�"�oʰ�]�l-���哻�|�9vcgV�h`l�+�
�l�c��<!)�8��3{����6<ǈ���������H�>�	��7���6嫉o;�l���:N,��p{p���/(�G�T�����O�׍y���X*�`���(��i�ъ\�/2��E�C^���B}M͒����6� ��r���C�<>�
���rup�	"�������h�IT��ymG$�q�r'vd��[j��.��-6����.�_�N��t�Gh���V%�~���!�Lx_�B��t���� \�a��蛠<�PX�%?����_��)8LM�9��U�����Y�6˶��J�Ę�i=��־~d��Ѝ��boX.�S�T�v`*ж��(&C�-n'O֧D:�����g�b���!��5��p�@.쿃aĮu�����j�=V!t8�SD-�T3������=u�v����M"5����4��l� �wJi�
P�tt�X��y�L"�8���y9��y���"0�"�
��{���@f��o��8d.Z�}epߠ�94�0��0w\���z��4�͞��lc��U_��g˒_^Q�R�!$~�/f��(=��׃�,{N�3!��DDC�%b�/���#���6z�b�7�V��K6%���a�&yR��!�	�M0�mu
��W���R��20�\ +룽���S0*e��L��:��>;�;�9�-�W�ǘ��]���Ձ@��޺���#(��T�M��oFb!�0�g+|���,K����])�6�3���@Q���/" ��:�z+��ٔ�DT*n�Lj6��4�O�P6i��i̖�!�p�i�"^m-?kȆ�2�X��W��y�4k�:&���Nv0,y� B���S�����O1T>����S�U�ߍ0��W�v)�<�H�i;5j����v>1Uvlq�2��@�2]v���~l�R,*AX���W9�H�܋�R"�D7��Y&�[V���`��Fe�]d]Ǒ�p���:���;�1��"k[��'3�Z�((����`�	��u��t?�Q40H��D�M%��U�ѭXK3��Ro��L�X�Nȇט�-W��,`���R��W�<�%�85YN��ow(m���iK�)@��-���6��1a�؏�d?O�3���x���]W�s�z�Cd���ᬡޯ�3�[~Q� ?�.�lyH6��N��U���zK��&gV@�P&�s��d�|�*H]䞤��0����pV���D���L3L����<����`��v@YZ
}P�@̳y�q��������e睼V!��!Y���B�ց�o��PC��>Y6���K�y�S���@����T��
�̕��=�VmK�F�m�2=	��s�;�+�G*P���)�fl�x�9�M��Zu����ӫu��a�*��;jobv=]���<A�-�Ӱ��7Wh��E�_Q������Coǚ��64N���ے�BF���!u{�?!f��d�)�7�64��]�\�<x��.*�w�������18B,UPs)�>� ���z1�����k�P
��`�B�7���ԕsX�ڋi�80�������+�Z�!?�K*��Pg�_D����j����g!�<u�ɛA  �y�)1���t�4��7�����)��ͻ�����&p��&+�o"a�iL���v��x�Ꮸ��bF���0�v��蜮�q��#���kA���;�xt�U����G�%G�ӂ���Mј�fB���Z��2����y]�"�f�Jc��{���臼�~���E*6����ʦ8vFm�t%9��>�Ď�a6!����Jde,��o%����Bz�F�	e����@��k���)�'�n^�8`��mM�GH. ({ὶ��pg�┩�Ƈ4��\�/�d􊄟|Z�͹t<rт�C�����7���@^&�-h&��"�>�F����g�E�[&%"�cv߰����T�K,��16�2<FD�O�H�(5(�m�t������zw�8�$����T���O����Y�����MȊO$���|r�����Ʊ�/�5PQ](�H<�u��?��f�u�<�:��"ƴ�/����Q>��F��sd��6p�M�j��ֈ�^x{�<iT� ������i�$P1	:�R<��0��g�#0�?�c�g�B�w���T�N�	yQ���&��ɬ�0�%�u�XsZ<�P-�pB�ۏ��p��b���jD��K":�����\��=I�2�:w��B�c�E�����U���N��"oS�=-�[Db����'e<6E�۟3m�>�V�6�*Ѥ؟I1��7���!�ʫ����2gČ`ǼS���"'S|����(]بvʬ����R��P}���偘M�uXf���Nk��2AU�@���_�H �[�������YI��[~6�����~�P�p�-t-�J���]�)8���-S���v+�6�&m�
��X�����@
f�R]O���⤀X�P�C�p6[�����n�t���J���M'��� 2�]ڵ A�痼�V6���:#������4�Z���eb���U�`l�E6? �3�<��q9��7�D�EE	�fewo��"��3��
���nv�,]���Br���"R��O�!��
�{��)Ֆ&�v�#`��Sm���4Bzćn��T�-@�|�½�=��]c�c�z�`(��D�Ie%G�'R�o�APq��.���0v��o�WvK�0�l5��B��R�<�kh��9�~�y2A��D�:�,쾿e�����٩9��e��������@"�w�7\u6f���
@�F�D�5�8��*$-�ug��1W)�}�9栆�о�Z��aV��*))`0�q�M	���F�w�ͭ����$�S���_��7L�h���K�z+�76v���w{��j�f~���%�%��&�Q��,�Hm#��l����� ��0>��!�H�d��pG
[�P�.M9d�ݩp����@[$r���䔵���4i��tK���@�p%�o�?�*C��>o��r�KW�S����K]��Ƙ-�L�fh�Pd�<*�_���a�ۨd͵�	p3�ݝ�b�8�=�a�rIm��;�Ow(_���Sb"^����0HdL��Y�0�Os�N/1o��<�V�G
N��Q�/�%��=%Ds\(rz����RwÄ�r�j��N;��@A�IG�H�d���A��UPK����E�;�ȁ�l|�.�FKv�dk'5V3��w�A�
vW?��պ+YBUso���F��H�l~�t�j\���_��c	˼I `��)5��Ҧ��>Q�J��TU�n�����S��b���Zb"9��4��'�d��zo���aQ\Yx��+��tC�{��Y�ɲ�=� ����c1o��D��2-�h[TEђZ�.=���=�����u����Xʴ�Y�0���P:�?2i5j4��?!��1|P4�[;�5*����D�
��H���+{�Kc���hS`�g�t�k��[Ds	��!��_|��$b3�����CWW�s�<�'+�-��^�����h!Z��X鎕ނR��m�e���L���[����Y�;CJ#���	cN�O�GA#��G�ɥBw1�lf�>SeV|�E��?�KB�X)g�l�d4��'
f��$����Q5�unZ�PXZY���b�}����O����$�$\��4Ew�E/P+�E��R�k���ߍi�u��ҺL��ia��\�/wzm���t̎"��
�Hb���W�oĵ��+!=8R�C#lX���>�r�"ܣE�$�`u���oSP"3�R����h���V��j����`�S�����@z�_s��Y����I����O����uaɳi��s�-��a�vZ�W�Β?�"�S���
 0�4F�_�&��1F�-�-�_������r̔1�'�I��(����gӼzN`Pk+�ԠzT#>��l��D�i��H��ɼ.��T	�?�1�-8zG���}O���ԡ���?�ڍ��e�\�"|{�ud�ߡ�]���k(+(��k���yoT�v
sѹ	�
�b
�*5����PD4S�LU�9�Z�1lq%�ʢE�Wt"r���-��p��N}�z�pJ)��t��I�T��
G*��z�D)������[��ft~� 3�-���2�`�o��J�\���h��Ǳ �D�s��U(�N������%yƎn��\�.��t�f��N�M�E&���nU���p�#j�^̒x��(;� �s���f�|p�$�j����aڸ1å��l,]�྄l� ��Jb��u��%;��H��rCi����Z����p��$�ߜg+�����Wف��"�T���|ə�Z������1���Y��� ���y��k�b{�b��<��MC(ԏo�����9G��_2$���)���d��t��;�ʤ��_��I��*�|�c�
B��U>�W��X��-n
`�7&:6�ћ�}#���fGd!��[�b`�F���,��K�G�L_���}�� ��>�:�<='8;��;:���4{AA��R(G�9�]�"�+�-h7�T��\#����	"�\+�t��]v)�uM��wɌ�#��]e����.�Q�^.`��1��>Zt"���t��������lѝ���J��JEme��,�QT�@�Ub������.A�w�c���X���D/��,W���켛r�66n�I��9�c�Fݟ��AW�tF���[��(ST�>�6�:�ҶC[-�2��}�ȉj�k`v��]�����(S�0n��+�=}ɶ	d�s�����2T��O(W(t�c�8�s�3<��%��{.0,E�%S-n���S�~Rf��gVy+A ��n'�mB�R����gX���I�YyFc
�!��A�"�,=�;�v۬f���P��W �����\3�mjh��+���q?	�/���,?��Y>��l�i� ��$S)���6I���e�/�)��6D\�j\J\"T�Tz Ch5Ry�,�fW���6�_�\�Eq�s�T�\{����XE\iI��E�j��99(��.8P|5�"ϾY��"�f-���)G��:��aa��dhW0�U���/���]�xE�=L&��&��a�f|^W��KC&5���]9���N�8GKV� t$�R����釘�EE�&k�? �;�� w�`����!�����������R{uy�W.��&�Ym��e���H����R��3���̆nB���AP����ep�ê��
�����q4><��^�a�|�{`#��woe���Y�X�rbw������4��I�A&�l�JW��]q���t,��"�D��*��52��w�XԚkR:1���1,1_��LJw
�b�As�����}��I��!�����4|]~}e(K�X������ÝmQ�(��\ �#Db'{���l����8���7i۸��y����4Ɨ�5Ѫ�[s2���G|�8&���������a'ʕ^ Y�T�:�:�6�I�0��/��TV���gu�]$QF�42cE�uxt�3�ӝ�������)Owa%.��>*��z��,��iB�b��6M���ų�+��Љ~w��p���F%s
d��;z���>��J�	 ��v�CWU-�_vs͏�X��4�i�]\{��-�W�*�>�s�����z>���Sc<8��9�k���ᎩH���2n�C*�fo�Kwq���cJ��c���\��V���H����hzY��sW��\v�0�-}���*�e�����e�l��W=�ԡˠA��Q�d�JY��Yr� 0=�½�U�5����q�+��FG�cs/�LgؼX� ����*`%�_�C4�q`���_FkD����C�NG�#�jכOߘCtA��偬{�ڃ���<Z�'�3�?�v#�eL5�����D9�Tc���P9/}#|��w9�TK���xXQ*|^��X^2��f�@]�/�A^�o>%<@�֊��f��&�����[�J8�:5�?�s ����xnw�}���7]Y��	?+'��a�t�K�YVF�S��*kN*��,*y�eɈ�G
lIӂ�`5�c;}���k'�\Ɔ.U���8�+м�1`W	P���jR{]%H�� ���ݑ�W) ���_�@��uOz��-Q����k��Go屮�T@��R�Pژf-z��E�B��ХjA��?�C�֓�@��Eb��ӎ��4�q8�g�bV�x����\UkI������^A�6m�tz�Z�)9;��HG��gM9�+@W�\��<��^C[?-"�ܝ�v���v�qs\�P�j�捍��D�H��>��J17�C��i�)3�g7Z�\|���c��	�RexuO��o�%}~�����Va}b�y�N��X�r���kT�r��	|��6F�ǔ+��7݄�Ĕ� ��
ځ5� �����b��'3g�L�do%�(����=��=DJ���ҘG�À�� �~~F�l�Z��P?l������eD���NI���hlC�������h������FA���LC��+�Ê��D7�q��>�X��W�~~���� 	���,��amO܎vѥp�l�3�<ئ@����:��7t/֗���S	qw�,KG�BpYke�su�("��2��H����$S��&�l���W��k���܄!h#�:��T 2�{8ߔ��
��
��Z�5��1�.v�vp����&f�0�����x��	u�,'ؤ�����ڐ39�䒩6wX��$`h?���#��@p�o9��$��+�RV��Ů6��Z��=fM
��B8~�jU����n���t5#S�_	{}}mxz�r�3NH�%��ZЩ�_\ ��g���T�LU[!��D���)�Dg�g�hq�7	�$(�^�� J��#־�	v��c�8���b��36�|����	L?���;B����)q�b�ن��$��4=�s�G�FM�V�(�o�g �lX�T�B��tf�ܺ�����b�#��'��`�I�B�&�Q�/����_�%?���X���MkT�g�tX����O�� �?��NL�#��&�<��J�Ig��OnXW+f�l�ܿ(�M%}_�)��A���0Q�B�$�M.��,�
��r7�g�+�-?�
�	(z���$��q(? ;o�]s8�c9�&D���=^��\�:)8#JY�#dx��;������M���A(�|�c��ʛ�R�o�&1�0��Ѐ!�.B v�x%dS��`�.������e����LBh���(�s�j�6h Gk���#JJ+Az����XGṒ�2�e����0.�U�Z�PY�`����f��W�3��g���Ɂ�k��[ӏ��]��q[OFrV�s�a@0��f	���i���Q���/���O��uyj0蘴����ö��G:����i�8g���ނ�,���" ���ю�����.<K�2u���c��pM?������ mr���O=��0a��8��'?X�!���:�.��94}4Q�1��l*�B���xչ#��	����5�!A5��uk��rp�S��Ѳ�O3r�Ϗ8rw�!�'C7����j��=?	�󗉈���f��S\��N.Pq�����?�T�\[�|; 	�� yW�F����枼`[����p�*ZyH��Mk�oز`�$���M���p�^w}��D=�������G�C���f��_���4�ͷ�|�����ځ�$r|Y�Q���S�F���t��t
��**��	ƾ�P4p��	�>���H_��/��]�ƻ�	A�^��JAb���oQ�\�t ��$��F3.#���*�j��[��-��0��� p'm�OI6K�Ud�����Y�>�7�hm?��2p%/0M������Z��êkU�w}��V�#����GC�(<$�r����*H.l���=Y������q�����0"S�]5/k��_�lVS�P�#k�'嬀y\��ڝ�n�1�������%0���E9�l�ܶ5����S΢u�%p\���Z]��%9�!-#^�!��j�Y5W6��K�K�q�m�Eɖ�����Pr����L�%*V?f:�5Y�3ܞ7����;}Hch�F �fr�O�	C�x�)�f�4�Ēp��B�b;�3)�FK��V_�deoo~Z��C�����/��߹`�ݓ�͋L*��/R��aN@�q�#��e^��r�we"���i��)Y�vq����G�>#R�����Qw)&�Ie������b�F��r�d��q`���>[��ʽ+�O)�ӿ��j���Os�.Zք]���~=:�OӨ��j�q�2�	���Ϯ4�U���L���v�ڙxƥj/�����-D,���=ׂ"k�0�%[��u%"���h��|1����'֌\՘�]}�lOd	�U<������*J�z�ؐ�����yĚ�^�s!��L�*�6��;����ЕN<3e1�#(S"�W��[&vçy�>Z�H(ܻ�����B���0-˘����97t�Ggd#�8���O�kh��[*W�,n�^ �7��"�/(1���Lnt��Y��F�*�Y���Ϸ4����G�]�"�3}y���zǨ慳A'Vp��AxkD� ^��˳��� �[�#LL�q��5����N�Z����2�ej?�;(���g��P5���@�Э�m��c���yM\Qk7Ե�XR w#�,N���7\H�ѵ��h[���Δ��FE�P�MB�X������)Q�q���~���p�pU|�>	���o
���a4y������������5z̠����U�ؠͽ"�E4��4l|�Wt_�v�^*F�Y�DnRe�C�����ȑq7X�4�����w����x��N��n� �Wk�k�"��Ƥ�5�n�
�kgv�#{wCcגܼI���F[�j�DF
XXN3PiE�.�l��ūu{��KU�:ut�G��#�RS#�����8��/����L0L������bX�S�]y����V�q�)��͒�D��FǍ[�5��f������Us��؂��z#�ӭ��L�����F�0�}������3ܥ��vA� ;?ڬ=A$�_�$0�3�[����^ߏ��T�O9.}��[o�!9�'�΁x�:(R#Ɓ���ꭔ�]���@笸���N�}Q�s̈�2��GB��-pT�BG��EcMl�?��
�IkY4���&�>���n�+Ȅ�B�b�/��ƠQ� �(�^�6O�EA���_=�&�b�v%*98����������1�}ǈ� .�4���Q��&V�SN$)3Ge,l��Y[��,�H?�٥��K��
BC+ͺ�ѻs.��4�6콯�E��:�iݝS��k������Z�`h�����f�eY�q5��(oU�
|�!.֗X��4�:�7ؾN2GU����?��������=�	��l�wR:�]��2�m���C����xR^E�#��EAt[�#�����<&"��L=����Î��o�=B9-�ޜ�fG�57ܵ�F�5-��07�v�.���sD��qH��6$�c`�c�� ��5� 7�W��<i�B�-ku��}s
fe�س��.Y�4׍��l�6�h�ߤ��� ��3߂��0�w1��ae��ᚎyg��8�%.R`,9:�;���d��0�w���~Ii/��+�(��<��A餞#�Ñً���E�]�$|EPL%l�4PaU\,�� �7�ҊE�?���+	���d�B�c�yE��鮏��Y�J|��y��������1��b.����T�,���1�r�(�(��T����Z���4;о	aʄ�mo=�3�W4&'��C��_�{�oS��N5��Am%��A;�R��"�o��+��H��G���m�i����Q�iC���vW��0���M��w�����ǒ��ڕ~w�#����er1�!�I&jnvI� ��컊$,m7.��G��@��l^t����~{W�شT�.e��њQ����:X�f/�"����`��.q��y�����ǟ�
/���k0Y�4{D/����Wd�@�xV����Y�|k�ߋ��Ss�=�,�������uT��yQ
좌�'���c�p�R5���~L�v������� 'n؎p?�9��ӻ���"�I?ܪ�Oό�v������2��$�l.M���v������:\�Y���*��E��{��r���O���D�V�(�K�"����8�d��j ��H����7/�KN6j*x��!�#s`�D�\�d��ǥ���T�avM�nA�t���u�a.~V�|�c��q����4��<�b����A�1�]��U�'�z �fx;Y�$ʆ�.+�E0V�xش����8�C�ی����~�����;���L=ǲ���UpMx���/V��,��s��S�.q��C���"F����L���&������׸�#�"N����y,w5�M�]�C�����k�[�&c�FL�*�m�s�_o�3[��g
�ҕ
��M������sC~�g*�����h���cv��hK ���%Tn�r&��[屚�yx�cn���ɋm�UQ��l���|���=�YQ/���ﶜ��X<����#ު���_�%MZ�J�\��O3��Ey)O�����V�0���w[Ы�!��������Z6KZ���T}zn�'C�)5�;��3{�X=FF��v�:C�R�����X`&s��8� ����� �����y������`l������/i�2W�@�Gb�0M�V�@���8��p���U�����^l#@�{�4�����5��򉵇�h�u{3��(i�,R*��^������)���2Õ��`Êe���i3*f&Q3=�)l��k���o�'�n��	��h#�T���7(�R��c�!dF��>�[�n�d>�X)�63�mơ8bo�|$y��	xMS}\�U���`7��C��c���3F���03�$�"%��i�f�q�u���\�z�������so(�p6�K$�h���ڌ�>��a�_Z.�T�1�xi�ۄ�I)&���D��2"A,~�}�F��K�	����uI$0�N>Hvi>��&�D4h��^�}�J�|���V_�Ǯ�z�:T�mq�@�Y?���P����Z�yMO	�#�g��lf���ѝ�����Wʔ���K��0�X>Ɉ���A�%c�Ó���S�X�8�x��������Ǚ&����`J�RN�u b	h�l�~�mFı��@�z'�AM���#�mvMsWs�G�~�n�arT9�,��-g��R���5�V�����܌G����z��TƼ�u���=D�܃���,PB�D���*�~�ʩ#�Mv8Y��8�?�k�޾!?Ԙ*v����8M^Df!xMPun���SN� "��a�{��{�����S�g��w�c�Y��v� O�-���H<m�F�}���ד�c!�~�!����&�M48��=@�K!=�OM�J�	ʆ �.S;�.���x��K�79~mqP�i:�!�#4����i�J�>� v��̓}�Gv?��Mѓg}Q�ãmݛ�ڥ ;[@6lƏM�nxAW���T� E�h���٠���:Li�uG�I�f�� ��.X��՚14�Cu����Q/�?�sk�S���;uf�'6�@Gq5g6���F�v)�Ix��TgśAV�X���m2�G"0�`I-v�'xެ�{��VQ���xR�^���s�8^SL�f\<�� ��s�2�ɨ0g�,����$�aAP1�	�y"&V7kK�_��
��eC'�Zn��e��d�����eD+�6U��|`�Z�r���A]T��x�.����v�&&�$�m4.��. ���w�p�S냔i^��A���Q��/���;̥��#��c�X�{�E�����
�{��n��Fq+l�&#�k�h:�-C�33t�t�Jf�\�'pKZ�����ϫ��Y���0ʶp�h�Y@Q���3�Б�d�7�d2�&`���W=ڙ�ܱ^���X�ߡ�ֲ �'�F�=��k�g�=��w��t͔� ��v7�79Oz��Z}�m�o�A?!@��0.����}��y�2�`8+��3�Q�G�C����7	��4�N.#!��?7^g�c�>M�E��(7o�-�ĔKm��^@�����������R�&{]+S���1�w�ɧ�8s����M�'
!xE[�1����0.���G�� �����[�JNq���d��'�:�y��w�`J�>��a�|9�ۋ�rAx�OB\S�H[�����m�@�X�ۂ��1'������>g��'-1+�X��+��Ԝ���p%nxB�'��a�p~�2��]�Z��V��|=�1��z����ˮ[@��B�0:��K>�H�n�m7�������4�S�]k����U���i�r[��-�c^�mAp�q�1�]�Q<�B�8�{���0��˰3|;Ύ��ߵ�6nY���LשwĐb*�b���V����a���2=Ӣ��t��['u�Lҗ8{!}����1�I�������
��]�SS쀟��eM�gٚ�q�/M��Oa�X�t����Q�>��Īt^JY�ExU#%�dgZu�]��܊(�ʀ���ym�馁gICI�;�." �~��y0��Ba1)v�&G�R0T��S��(ö�^ȵ�-�ayF{�R}���-�ȼ�����~�-	.c^��lxŽ�E�IY���Iy�N~Ch��5|������̶T:��CC�eM�[4�5�0\��g	E>ߎi�}��ہ�8���#�mN��z�Z�I�0���Ի����w_��i�q��l:<�׍��v+:��]��_jq��<N㞋��}�����e�d ��<���[��>�J=I�e�ơ=�&����Z� G"_�ͬ��C6$��Mp�+��V^>&��J����p�bK�u>R�%�B�������:�[�C��ݧp���/]'��m��\-;�c�M&<�}œ)R�6���]�}�@�a�\�R��5b��T�v����.�ԸX����Eڅ,ɀj�'�5lI+tڍ9�6/�=�4���t��#P�q�}�&�B�GZ����|@Q�.̓%�DͷgDY�x[��zƶ��Ne�a�D)���y.=���&B�!5���*��yx}�1��M��C��߯8�u�b��D��}|��$&���b���7P�Q<xr��z�V*�����b=�����.&=c�M�� ���m�m�(����(Ų�4��DC��Y��>�-�7����K�%;M�u���െ���N�Vo ���~z�����7i�>43�2H J"�"��0���R��,��;�fxk1��`�����k��Ducď���׳׃��Ї�������,��7�|hL؅�#�H⼳y�%!�ٵ?�)RS�@j�"~�G�	G}G��>;��;����y�	��1��g��d�?i����s��V�`�iڟ|*�\���r{�q:�;�Nwo�,��rPLFא�<	ro����ǚ��1��a��>�_k��@෠�3U���/��n��~��9�3Kq�=o@'�r�*�Ӗ�r��mLØ]�br�t�2�&���b@�u�.〕87�šH�m��%lT�3��O��j��9͊V@ �
�����1��2 EEjQ���=��4�
���
�LJ�����!~�i��8�Ñ���Ʋw������ҙ�;YJ�:m����o^C�<��������D�а�"	֊���21L��J���'��{�A~���mj-��~����!~>���!�	Θ.Iiǉ�b�2�&�g6o�#���,��@p��������5���g�O$��M�tR 45�E���)г?[A�v�1l]��XG\��"�
��'�%՝R#%:��n����ᷭ1^�;G5��M
�:~��b�嘤�K���X6q����
��[�@�oV�k�X[P-��m�X���u��$�j�g>���L+[o_�,�)���H)6�υ$�����6�?E�Gq�"�A�kV}O�c}���"$¥j��k�œ�K>��6�,p6�骀�AZ���|Pa�L�@����A	V0�����`�/����A
& �vK�C�6г3�)��s
x���*��� �t�k$�d2d�L�O�nqD�����,�������Ryx�+mU���=㤭�k���
%����o�ӵ�OZ�!�n�_I���h^��LG���f(*�mc0�jT�7Gwq�#4�n���5�pt<�����VS\9�,��Bb�`��6Ne�T,"�v{��hlF~#�GY�m�����*�{���T�=.�E�T%ԋ�ZSm*[���7c�;ag@�3"�L��\կ�l<�Iz�yR�Ia+�i��� ��5�z�\�3v2�G���xv��6>4��g-1'��)>�HI֚E�?�`�Ђ�r�m�[�tk/T�6���L/��N,K��.S'2�:ϑe3kF�CԠ�?�f���h��n+�u�h?�N������8k���H����"����d�}���Xo�DN�06��Rddx$ݫ���� }&�b����TI��<�J��-�ׄ��|よ-�^A6���ID�N�1a�2?�n��߂�;d�N�ơe0�Æ1�+��ێ,���爵�q���L��3���LPtf��*��=g���U����쥰{*f�c�8��(ʜ �������D=�}���#Ro?��H��g�*C��lQ��4>bnL�L��G�b C�z���c2���c�:"}��L{�ĸ�(�pz�������@�e-�]�+�,���L!�w�����`4����!�Z[I@�I��c�7�6G�*��xF0�m�NZɃn���7��˰�+r���<((����4Y"�j�i$z�BR�J���Z�p�8S���Ȱ��!v<L�n��2�t���'�ݗfjIg&���yi A�!�wH�曶2�n��`^��(�Dqw�����.�D�#�gTE�E|P�@&���*R���}�;0no9���d�A&\4�h��h��II�T#����m�'��q�k��/�@�}�f��E!NѺE�|A�!l]_��e�-�5��86 �"f�_���f��.ש�����g)ַʫ4O�����Q���x1�OM�z�ɢDL5�9),�!IK�<5��B�&պ�i'�8��b���5��YI*�tʦ��y1����S����s�!�b���V0����O>��C��a#<eΜm�s5������D�fQta���8�(z�����5���5'�jK�dr��=C4r���I�5��|l���Ҙv[�'���r��[�����x6[\�kPX��]���-jL���ʆo�&ݗ�R��n�a�u�4A��2�PEXtw
Q���u�TF��E�����4½o� +8�_�kUi�V��e��K�d�ى��%����}�	O�ן��B�K�XfD���P)���]t¶��FT�\ ���5ݺ��!�r��rZ��ռ뾹��sX�&��+�T��t���3���D
K.���]d� U~;��N�E'!�@�/��[�������� \��@Kf��Ey�*���`.��6�m�FDJWe�,����R���)|t2���H�5�%@b<�Q5_�P�	�M��^_�B����v�#�6�7�[���y�S`Z����!ɎkK^�N� ;�Qia �/F���ŉR,�G����z�Ѵ�P���ˎN�T�W���Inb�}NS3��`Ӧ�S&as�6\a�7�Bw�̤V�A����� �#�=��5؏0L�t�L��#�x�w��C��O��yK�]�,T괅���iD���@B�w�0�=%? ��C���^����H�F�i=��o�^'�3Jh��AG�G䇍Ϳ�W��f�@���C8-hj/��_��� �p�B�,$gP�����A���x?�_U���.�@�G^�@)��}<�.���<D�����Q�:p��ϥ��XLϊ�V�|Yf?\��V�ӻ�_m�^7`h]��9 �A}q�	� �Ӌ&jR.�bwG��5z@%�)��)tm��xz$A������ Ȇ�^�1�%��Ѝ3��ӦW��2+k.�u��:���\�eD��g�_x���2Z@J��eQ��q;Z�6Ҽ�6��6�"��3���ޑ)ʩ`��e���.�ro�87��#��	��d�UB^h��D���_m��34Z�g�D�S�X(yi��{�%� �&��}cz�T�^f���o�wa���>�X�����F/_�| �Clt���@�^�PK�|e��Xl3�xG�\�b5*ܷ�~+1�.��m\���k���*R�E���(ˋJNPO>�v�7���T�&�Q��\�*r�qZ����p{�^l���E`mӤ_����۠����$�2T��1�#Oޱ�V-Ŝ�ԝ�^~5�+�O9;=e��s��c�ĥ@}8y{L�ӿ� CJI$q���K�s��tt.���ހ�*�M��ge+D���`T�0��yrg�T
s�a}��q�שDbwA,����n�����N��� �4�H��R�ㄞ-����&}r�"�����m�U�8K(��:�ؤ_B'VZ�v�q�2H-�^�������Y��	Qn@�2��[��M�����L���@;B���7�Y���v�<v��v���~�jZ�T2���z�����j���t)���E���_e����ޅ�|'�m�An�k�J���A�R���&Y�2f��Rي���̕�f(�Y���>��߱������:A`�c4h�~��tb�K_�F�MZ����&���u����!�HW%t�Q;����ef������ 4JiH^=�a�#N��wH����`�B�D˯B�4�̇4bB�'��ϋ�X�#�[�jt�3�=~7^�#����!z���9[؝dY�L��y�>�g C���x՘*c�=�Hf��٪^��
HHUj��~�[tD� e]?��`����a�V�.�t����p�f��w�
�6�=����p߸�j�}O�:�j&�����t���>��({��n�����G��C!uz���j)�d}��[��˩��ۤ�b�Ic����P��ok��1��Ύ�_N��y�~�X�2Vh�ܧX��a��exо�����at$B�r ����AP �s�f���\���a�#y0��I���CM�ac�["�[�Mr���`���ۊ��f���J��� :�L����خR�l��*�^����-j4�2�фF��~F���;��Cž>�Kee
^�v�b��,yT����r4�oց��5��SpAsćI���������@�t`�E��E���Ev*��5l�~Yrj��O-�/�Ӻ��$+e����4�Ҵ��=1�Y��Cxv���`d��~OV���c!ys�Z�uㆊ!vIl�Ne3��mA�HrAG:�v ��r����z�t*���1!�j��_d��y6��4�n�;�Q񛥩��a�;�q�P|�~?x���I�c�㿲.L��Z܇�Y墻yi֢޸;�B�&���� n*��wFlѨg�ߞM
��%J-Q׆YUK��܈{�?s�'���$��ݨ~�X�D=N7C<��K�<FC/�D& u�3���%Q&�;}��tO���#�æC۳��F�8Я;)���|qi���6�Ie����g\!���d_~��C; \c�x��X���#KM��G�S�
#��g3�喚���p:�QN(�t�1�S����O��~y��TW/0�.�#5"��Up(��~{���G���m�^��F �)�6�_�I�OS���0�Ɗg�k�nH���Q��Rl\i6��@H������,Ӭ|J�R+`�n9����F?��$�Dh� �y��85F��������I5Nx�!@��Ѡ)L�Yt,�j�E@�K�y���	�ɤ�k�a�ѢN|�����O!���&:��IO�X�[�BN;
^2٣D�y$�.ؤ���i����ߔRZ��lX�n���q��� ��V�TR��V��k}�������=X�r�����Ǉ���/�o�''�:ؓD>�~*�-^�p��n/ؙ�ΑJ�.���#�����X���A~-�-zѬ0�$�̿��x��pM
]���a=���_�o 6�"�Rx\W�J��Es�k�C�',d����X+ay*z��b�Q/M\-Y羻h�)H��K�7J����r��2r��ެ�&O�}�c�,u��6�4
\��`Ǚzzt|�*Q�t�@[i��Q9�G�z-�/��GݙX;|P���(��A �>����`D�k�h%�%�?1�RfC�kS�P6���+�c@Z|�|XY±���eyV�뿱g�g���<�]룚��7?#1u�?`MNo+RH4��s+vp��=��`F�䰓'Ō�^�Qu�����!��Yd�@9-�P�b�vZ����Wsaa�#��Y:�gS��Cp_@���-����#L���|��B�4V�ԛ�괬j�	�юԶ�?��͐)�g)�h����#E��_�� /?�.��l��,�����j��wQ}'Vr%�:8�
J���>�K­{'����F��"pxn�K��2Zg �@�=�©/�"�Wv�
̤ ��2���}o��<��y�K0�ʶp_[�آnk�5H�&�F�j�%�41���c8}���ǩ~$��'�����[<4]���j�J���m�(��(Ɗ-���E�ޒ�c�aB�D����|�E�e��0���H������)�-(q-�}r���R�z��T�(���i�y��	d(*��H8��b7ԗ���z�|Z;p�U�6}����H��Ó��7���)��&����T��&�-�DX aط��:ʫ9�jz�|�P0J��~f:����ǨA
1m}�3z3�����F�s�����.��j���tв��(�ł%�a����YR�!q�#�"�X�gַ�9��_�>�r\�����%��j�䷖�,��<�P�d����QT�N�Dku'\�>ɳ����3~��e�D4��гO��2gd�?�l@I��Ԟa�VT^�KLXbdE� ƮN�;�N �v{�	�]�����m�N�t����^I��w�����g�0b��X��}���󶩀�I`��Z�Ni�f̤�ʚuz|(�հjhn�kh]X��E%
��*�;�����$���ʝ���L9�wId�=��TM�����9*~�Wk\%�a� l�N�a�	v��?K[ق\������k���D; �-��Ǳ!�w��2%������&j53�;�O�x��.� : �諴�>����`8zPZ�0Sْ����rD�s1={=�i_�%6���4E��璎j�����}��ǃa�j�c>m�3w7���X�Z�*xPS��h��68�<�ǡj��&��./#�D�&���ZN��c#�k"R� �D�P3��!��B�`��4���r�vymq�w�YMn�{��X5lp�&=&c��q����@���Bg�g��d���2��B]�������^p������Q������BN�E"���e��9rY�((aV"E�!4����K�QJe��ȀHe	��	~t����Ⱥ�Ѩ�I�
�D��:�!��h����~T��5H,�4h.�$P�����Cc ���-LH���el�f��jh�d�B�/��#!|�҆��yFι$�w��j�1��j3S�)�Y7v������l�۔2d���A���wԉ����
W�����,�>C�g���"O��ݍ^�%1V�S�\�`6T��M�چ�n�o|�H��%�q_�A�б��������sm�Z�m���>b�W���g2��𢡊�q ����c�G�[{��"��D�<J�}�o�&��cΒe�e׽?w���"W1�S����#v�9�ē�E�#��@i�K,B���I"ޞ���2������V�������XA�dR5��B���jV�VLūCO�H=]��<���#kbw9HI�]�<�����E�oo��5�v���#�A��j�������N����&J�w�u��$^0��M/pk�RS&���b��I�R�~�.n'�2S`��,�H�pqf��}ϭc���Gҝ��%,�P����
s��3��(�%�}Hp&��{H� �!Z6�Iү����I$i�Iü�KP8jc,dćR+5CL���?��Q���.����?�@������9���Uz���3S�W�a����(�v�������������PSZ8��K\����e׸8t�G~��~d����I _m�vF8y�.<Tk#�?黬mvnγ��z����v͜ )j	�Gȅ4τQZbK�!yY��󩺮;���(�t�LZ=�nJSizUKb·2��c����LL������\˕���
y�mp�M���~��I�D�0�c�C}�FQ˗��jJ�ɾ~���!�P˼u��(�Q�"Lw_�^���]�䚦�����T�xRB�z ���є6��%d�ɣ�!*��t�q|� ��毤M2��|��Df�L�n����]��p�鯲�	�g������V��z�E��x�n���5�����Q��4�F�:��Y�ϧ�U�a � ���jU�';'�l��|T��P�J��\�9����$�[Y
�M��S��ۥ��f�!íWb��
��T�-����|�0;܆b�&ٛA�m}�2�r��岟H4�gݹQ2H�y�sZ��|��۸>-�`�Z����IuT��@;��$�Qѻ�? b��|��@�^�$��í�3�ư*?3�,8� �5�6^�?�U�{�޷X����Sm����bM���2F��;F �����B���?�m5ƿj���E*�h���(�P]�)��k����w���#����C�?�Q<��F�"ԓ^�@Z�O �U��:&�>��~��`5���iB�ë�����h�][����P@������W�F0��g��|��Ɖ��I��Y/rxF����Ƞ��G�VY4���ֺ˲45C�9S2i	�m�Y����&�g5,5��m#S#
�	��|ߝ����r�}���1$a��k�;�7%Ļ��w��A��8[R�>���Z�K݀G���T�GI �!�x�\�ttH5��yL��l�N��nK���]PS��P�|
|���8��c2lS���ɦ)u`�x�0�̌�V��J�e$�ð#���#�����}���`�zAe0̙<v��>�F�M���UTm���3������f@�'D��9�o��$�nat$����Cȣ�i���:i�V��"G���D�Pആ�愫����3����%%G	���%~��l�95�9(⧊�+�^�ZZفפ��/��߲�Z&a�zh�.��t��S����Na?��{��Q�=w#�p�Ŀ&|�k)�ЄI�t��2.r�u�6��h\%���te�]⒆��3�B��_y�W�Ʀ%�I��������!���L�)J�fs��5���@8N/].)��Fz�|��É�l�q�Ω)��s��C$��Q|	c�jE(Z[��G���[��/[߻Ա�I��S�xtD6X7�,���;9W$^ZX�ʑ<"sU�n�	��"����Q��T��Jo��望͆=��vK�׺��5�3��(-�i��ʝ��N��C�%�!�.W#�H
�,�<s]�;$�@&:�iwJm"lks
�N�u�&��r�S����XQ!&r|�g���*s;�!-v����B�U��wu��Gf�~E�	��odVQ��J%j�y(�)�C;O
�h" �?i�x��ױ�MZ��`B�w5B�xeÕ@Z^BLS���̯�,������}K3�n`IUz�g��'c_���������q��orْ���oq*r\��Miai2��5²B�Y����	�t~�+<R]� ��i��Y|�Pޟ�_�fG0�;6y��gŚW��
0Z3��z �E�w��>�~�����EeI��z���u��z�zPD+P���x���Y&�IwV+�/���$� R$u�H��@�罈	�2��E�r��7M�ر:%$5ʹLȺ�H�U�����>���@��z�%�,.�2oF�0���n�S��c�1�N����!���B��-��r\!ق⢀<%B`<W�0Y.ֆ!j�c��|V}��X?%w��b��dZ��u�k����J4���z	�`��E�!i/z�dZ�i\S~�OH8,�ZfY8�v4���`J��1A�����hBl4�q_�ȩԼ�{�8~�8�������uy~���@,����a3���xnF�h�<�� ���q���0�K�6N���Ve����]
�E�d�W�M�x!`>����_0��](�B��B��S�C���5�aX�Q�ߍ������w ��Fՙ6�J��2����{�N�ͬC䝌�KK�ޤ�/L�뤡l)��7��>9Fv2ʄi����c��0�u�P|7���٫:(�F��/�t��X\SS�$%�
�V�`��%{iV�6l�o�9T{{�O(���� t!��`n�toV�>�֙=&Dbj)|�I�Y����!s.RT�-V5��I���{���;xJ_sR�Mۆ��$t��md��m0���W�y��� �Ǌ;���0���0l/ërkT�V����2Lmt�.nj8D0�◶�����*�_�T͋h��w�;�>����d���nZ�
�pͧ7��������!:�^BH�`$8��_��nk�4�!�h�RD��1���CFO��۠���𒝖e�c�MvUA��Q1?�2�� Io�k�1d�
a��R<���a��7(��D�p���%V<�2��{*�(��ǁ�s/L��������G����1!�`s����@7�9Hf�z���ʄ��އ�i��
K�5�%���g�nJ�R#U{gb�`���J��v>(�4{(fӎ_t�!����Ã�"*�S�^8���b�mt�; �w-���@Z��_����I�S$������vuX�un�66W��F��(i�ȕI���V��E�$��*c\��$�-�\ s�1��ȝ�E�Q�y[�&v|M_�=P2�e�~�����Pہ�7��p ī����`��		@�G��f˴qa�ԇiD�҈��Cw���[{����J��s/Ĺ/?@����v����#��XWr#�<ؘ�.46�J�����A��a3�0t�PX;�cS�Ӫ��&+_V�ٵzAp��H�VED��ɋ��s��y㐖P�ۃ�8��vf-7or**�{{>{��u�~�:���p���I��L��<�d��S��䁕�į�����Q��9\�H3�o[m�m
�
�%('�oh&	�{����#���r�| `V~A�Ra�S��H �%�pl]s���?&���Ir*�$���\�M��V&l�I���-V�Ǐ��7��6y߅\���0qz53�A� ���<�Jk9�����J��Bbe	I�ƽ���骴 %���ǒ��=t��pR �������V�p��!�&�G��T=�FתH��0����ŎD~jB�HR�0M�|���@��Xˍ�� ��߄q�rR���A�b7�׉쯋�b�`����J����~fn�h�-�9���u�v�{�Nk���p���9tL�E�e�ڏ��GM�oT���3����s+mA!6\���֯�!CB�V:֏�j��
�7��@]�{hw`���N�T|(�Aa�����F��G�~Q)�`ڟ~�>�P#�ctlo&P���ml�w3JU&�j\��уH�ԯ��ck��T~��rTi���$��h�xP����Z�jW����K�Yzc��^���Vm�!ǂY�����D��|���ᒱ�@�"���3�{�����۝�C29@�m��)��&9^I���ǀ������ۇ<Zˉ�~��]�i ����l���o���ɘ� `�ؓ:�CզA�:�VUt�K������~�]���7��p�5�U���턓#V��,��;�' �^�.��Dz����`+����	hK�N�k��Y�}ؿ����p#��EMvߞ6�fӫ��p���IG��KZ�T<��AR��3k�ø����#�̡�c�^�+�n"D3���e�
<cl��\ ���
ܰ�d}� �oڇ��jl��à����X�-�
\�[�����yFR�J d�@�߲�֡g�LZv Uk���b��8�k19`A��ˇٌZ�LRj�=�"Z�8�$�дr����]��\�45�w��ئOa��V;��M��
Sm�,R%���Y��V���)Shԯ �2�#xϕ
g��u��5�bR ��c}'���5V����_7c�<������w�+dV�92lg�?/0b��-h`��u�X��
�2�?E��|L�10�qٻԶ
R�RE�n�̫Q�C�����Ym�;�)�!4,;p�K�����4}	���"�_fc���lO��R@��c��^XHP�_���'��bgƂD^�G;Pi��BK����o���P�n��"&0?�"�k[�S)��<(�QW ���LN7A�˰�ΰ�D�B��"?��bOy�\�k泦
�P=���Y�t=YOs��p�>�0�����Ѯ�U��滙Z���`P��"�)ʓ�<Q��y�w}JV�6�.�xi��:Z?$�k,w�0�47�����>���X�xkN�Lp�9�ҿ��z�F˹0�S���~��ڮ�1��g����s���"�<�\�zD���v��Z2&\ZC�v��#X�K�����gK�3��b��&N)1�!&�=��͕�/��b�<�im�[�Aߥ�md�ܗ���T8�)lO6�[@n���54�l���)~G�g�o�X�_�'�m
�v�݈]A4˛䪊�M��Gwa�>~L��|���0����=��E��t8 �tҮ�N����^��I�r��c��5��0�*mK,�`���1�͠��jqp?������v�ӱ�S6LI<�����6���`|��s���,����M���mH�����u��m�u�<'M�g��r��v��=!���1\hu�?7��R,���/�R�X�ru�])oe��a��*�n�)c��ި��k|)}�C]��<b�U,�RB%��I!4�i���_/�ā�VG�d�E�f5��i+��@��dɬ[��������ƕSX>T#L�-��G.��A��Y�>>Qy�Q{"��/�۳��!>Z.�b�>[A���t���ݲZ�!�'C."t�k�=I>�z՛F��HV���rc��8F��9�il�*����h���Q�L�����<kK��E��l�Ff���<�h�JO�*�K��Л7��V�GN��4���8|z6)���J�%e>=�v�5n��^�uDb�
��k�	�;����6#�'U3���տ-�~3��%D�Ű��CÇ�ik�*��W�9�>?��~�b��VO�.֚8�6���JcŃ���0���r��\�	�vm@�c��Ӗ���	���Lh���$�B�\M8(���?��'���/ﬔ���N�@��{E���w�!�T��tX��PZk�qDq�vC:+S��O|�MK)�8Z��T) �|՘�a��r��LY3���܁����E�2�+�j��E�6�a����w3�����>�HP~9s�E��4�Ψ����m�$�촳Y��=R��˦ᠨZ�J��Hxl�.2�����lI�"��v:J�����Q=�Hg��B���.�:s̽�s���1� !�Wt��J���?c	=�N������ǘ�u���B��ދ+"e !���"l�~Zj�Ŷ˱�RN����R"'�4f�Ë%�z���4��Q�8t�6Sd�r���hM7r+Y��0�CU�W�������p���N���e�m���\����a���q��Ғ�*� L��K^��fk�-�l�T$8?��Uv��`�R�:I�s�� >�*��\�en`�T�Vd���c{Q��v_V��YK�X؝�g��OzH��%���h֝�iO��{J����y<��oНJY6�u��1��r�3(u���k!f7*�/2PA�6�b]�~Љ�E�qG\d�Ŕa	�T���[��Ri���m�P�=��X/����w~���s��x!�����9���C+J�����{�h%,g��^;{ݽ��cH R����c֕�CB�dO�ى</(��P��&e��t���0�r� iPY8��#N�84o�����^F�-��*
��D������ي�,�X̠U��W��	`i���t)J����ھɤظ����p��44~SiE�4�]�Y����<;a$X��Yua��wȂs;lrR�׽ �/������`;E����p%t����R�pu���%���X����;
g�:j]�a;�D�����'��] �[a��R�p�=�7� i�y�Cw�n�pL�[z�
еB�2)�W�@;�#@�r�}�H��'����^����1�˯G�|>�B+e�?ƫo�3���Sմ)� ��<��"�FAa����z��.�%_3�t��ǣ�2ᳯ��H������ϕp~�0��K�&�,m�U����;��r��<�� ģ��*�>�V���f1�a@cX:�e�����bB � �қh�IO����<��4 �T�?O��� {�YJ�������lD�=O�wl8� ��%M7r�i�Q�P��a,>XW�N��k�M�/��<K��͝4k���e���S��R�w��]���O ,� >�t���gga ^�-\�D@�kb�]��Uψ���U�Dh�~D���1���`##�g��o/E�8���,*˕��k�L(��ίior\Ο�|x�}`r1^�Ē��\6ֳ��f,�L�.�~��\���꿸A �]Ű�|x���B��8,��x�^L���F�O�^���N'x�!2����K��S�5��ڼS�Ƣ�E��J�vm��ͭ^��-�f�9�ҭ���ñ I�)5%M*�n9�U%�v_)�F�m�WV��H$�'!���Ⱦ�"4�
J��n&�e�h;nYPEo����YC��b�A��"F�?Nv�~η���L��6v�	�n���&��a^�
[�l�Z�=SIq#���UO:�C�����F�ƻ0���"�s6�r
�`t�.�SD:�aٜ��a_�N���������~�dJ�"�re�^~6�/�%!�V�y�Ӥ3��g�@��Y�c(z2�p�+�K���i��r���Q���f�1am�B/�6<��+O��?� �^�=���� �L|�D��
��L�Z�Ww,�Db�p�Yq6������j���hS��d[)i���3���#8� $.U:^��#�3x����W��V��3ːύ���r;,:����[�O�~Ҕ�Fu�3�ڷ��uz8#h<HY�U"
\ڤRY�֑�%2�7�1i�6qo������""�<�8���e��-��#�����]�=�P�L�(�[1N;��jI�8|H��M��J��͠?G�B�B��:�BCq�g��c�R.Ɏ�z./
�W���na�D��W'�c��,�X��c��nA�Ɍ�1(�;ׂ�\ge�r <ޣ}���Ҥ<�� ��s�";���7�y&W�{�p��ʁ� lu�zJ!/��ރ%��Ĺ� ��uB)R�@@��4y�Ek�
u<�}+�@���١c�Y(�Zz���~���ӧS�2Z�AcNZZ�\m?�'��[T�Ѿ���q�O�`�e�W���ĝb����^�KK�����lX����B\�Ծɿ��Eķ4Z�\%����M��!��#'@�b%CEL{�~c����Ý��)d_Z�ϫ�C\�Rw �)�s3~�'�[m25�٦(�W�ޭ��nFz@"\πFP��&]��I\��LM�.�)�o�_?LB(0��g)<�Ƅ6L�Tė��ڋ#}a�e+���DziK�H�wd�t�BｦH��>�(��g��xy'z��vSoD�\Y���8=�`�o@�-���.�m�B�����J��ݥ_3��m��i��*;�\q��_�U�3�dO�A� o]ˎ��!�Ƿ��)@>Y~�\_�޷�i7L��h����*�JsH|ʋ�����"�
0mY������%ی_{��{U��ͤ��;
Ӥ̤�k��:�&as:}��z?ߝ��x�sQ�Ȧ�t�332�VH^��x'¸�.�c��� }�Z�g�^�	]9s�c���T�`.lEh�n��w�m�.���&��ʊk]܎Mj-I
���Q��Y��
d���  Ĉ�?�JM�"�$� ��q���������m�k3����n�fR��cb�{jk��z�5nڡ=�������U��%���o!}���i�ט�J�jf�YXnۛ{��'-j&�����\����S���VF7R��T#!�6yt?��bѬ��	�q0
%Z�P�CHy���;�tc���6�n|�巸���j9^��LצYx<fIZ���:���7;�<`�1�ڴ�y/��p�|'Oh�����8�*@fl(@��d��9�\V�(�|RՊھ�2�"�a
 0�AMj�+�p�bh�0��.k��|$gCl�,�2c ��n�:��Nݯ�T@�W��H�av	��X�a��"	�a*Ŕhc�̒%%�^
M�Õz��]�EI���;n�����O:LlO��jD8\	���������p�J�e~_rqv���>m�c��z�%NzB�\-?�T�e2�
:�"�)�b]|:�P�x��R���|�������"�βXլQ�?��jy7���H�X,������&J$��z!�!6%F�T 8�N�p�H� ��cE�S���Fܐ�	xQ�s� @L�W�$T���O����P�BEvͬBkB��.��h|p��s{g��d�;m:���P���`��X�]�k|x�������#n���v�Z�����M��d����@�o���g|ى��Qby�dN]����Nw̓���(��X0��&6�$IGNLA/�b���ÚA�?u{��&?��_OAD%�9`�T���Uҩ�We�R#02;E���\dU���L�	sj&Lp��vM2�IYB�����O9�q�gs{�U����P��ʛP�\�64ee(v��[%�s࿠ѧc��N����]�8&ۯ��P~V8�����ݍt77����W�D�Z��(Y��͛�q]Z�R)�YZ����Kj��G'r>����R�7�~%��<�\+����t�!<�)>{���j6f](| ]�m�K���-{ |@�dOv-tvH��vٸ:xU���U7��a��ec�^ވ��=LF`��	�(�1:�@gB���v!��6#�W�\���D�Ǵ��O�@�o���V�����zRG7��5�/��������ԓ���MMG��o��[��+I�������߬V֓�=�"�f��C`NJ{���(��A��o��`�IZ4��ߝ_�Zn1�خY����D`����ʓ���U)T�LDx�KE�:(�o�{�8*s�z</��Ug���.��sq����\��B>~����L�!LC�ʁ�ɸL�b}��a0P#sh��-���ĴK�?&��Xl(u@ R��+�L�p�[����G{{AB1���,��)P@P��Sh:L���g�+-Rr���!�w+ke��������k�^g�<��6Ħ��2V������TV`X{�`�
Lh���EэP�kA̋K�6��6��x��Y�yV�����'Eו���!�І)��ӭ���;��W�������ˈX"�ɤu�`�}���P�x��ll���71c���r�#*@�O�.̖��[�d��Ec�N���ݱRb��M������@h���+ҹ��ԖݟA�4&�u�4��ˬʤ(�/�Z�	��,z�G�xz�JԮ1�t{�Hz,0��q����.Go lC�$ui��՗^����恗6l��o���AT��<�C�o�H@j����$<�3 dZ�Ԭ���8(T��⃎{��kqzx``��K�ܠ��.��u�jB�{�)�Y=����
^e�:'��{�M��1u~ޯ��>#�৆G���T�{r��Ґ&����S���D��eE]0������[�*�\�~Gϥ�6�/�YM1�V�x0�ҚP�*zl�t��G
,r}�-�S�jhߢ��Aֺ���#�cz���g*��6ku,��@H������2�:�X�"�ۚ�R ^�L�������������������#='%�-/-#%'%#=?=#%'$#,/-#'%�]_]cegecmomcegdct{}c-gec�mc�eec]_]#%'%#-/-#%'%#�=	#%'s#~/r#s'`#�ߎ��������������P��������#�#%#-/,#�#%#*?=#%'%#)/-#''%#]_]cegecmomc�fec|.cgcocg#c4_1#@'l#C/K#J'%#�>=#$'#/#'#�߿��������������������߸#%'%#`/D#F'W#R?N#J'C#Y/#f'J#/_-c
gcocg
c}cSgnclo+cg	c8_#@'W#^/D#J'K#=?=#'	#/#'	#������������e�������������ߤ#W'L#J/E#Q'%#�?#h'L#N/_#J'V#2_;cgEc.ocgccgcocgKc}_#I'I#/_#L'B#U?I#V'#_/H#V'@#�߫��������������������߼#H'@#-/-#h'L#^?O#J'V#B/K#Q'�#}_
cgc	ocgc�]c*gcocgc4_3#B'#~/T#V'Q#X?P#%'%#/&#$'u#�߲����������������������#'	#/#'#=?=#a'%#,/{#D'W#_4c	g c$ocg
c}}cAgacmo9cgc3_.#I'D#Y/D#J'K#=?=#%#�'-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������H�-d,8�ECp�*����a�������MU�Q�=
��~�mӞ�!�����8V���'����i�=l�Y�d��z�����y�A���NC��6����aĎ����r���/�W��زs�L%0���N8�&��l���K֞�����tsU����z�
���FY��<ܷ�!�pɺ������#�n�*��^lkTB��Ğ�H�#��M�V�8s�t�褂��=��� }"oߐ�����@5�C�)����+��oBoh .�w=��� Ł>p��:&LP�w���=N	�:��'���6ôx��Z�������� ���R�.1C����"��s���+�\�Qw|j����@����y�p��c:*V��il~�}�5��'����>K���^P�#�@	��qW���d�&�C��P��k|;��?Ԭ�s�}VN�PD���?(�rG��O¬i�#&�����N�����C]�*t��b\|оa�ӷ_��=�T����޻neU�ԃ��f�'@~���B�f^l����&��Ѻ��
���*d)¬+���Y҈fE;��2Lg�/�fElR��pPr�ٌ��DOQ�.UI
�~3q���(�jj�uiN��Z�G�p��(�����#h��پ�����	�~`D��dFB����3JF�"�a�}Ɋ�� ���1JI�Ś�`������O�ä�b��`` M��O�2�����ԥs����b]@X��-�A�k*�|����vɛڶ�w(����xP+��wW�0�����_�km���._:��JVn� {zHLd4t��m�RN9$?_��Z����A�X�.��r�)�S��J�cp@֜fW����;�e*C�a���D�/�db���JP@E��J��O�og����JaR�ޔ
L��ދ�w��?���c$u���"k��[�*�T攳������ƕ����0�ch��w!$��H�,J(2�K��Ps�y��8�k"�46Q���
����=
��k�]�0��{ty,KW�-������
c��GY��jk���F
�x���[bi��>�p.��FH��"��Na�w�}D!�$�|D���T]�m��a�5m�wX�a��U�le�Q�a�m$꽕<-̠GL�{�+�!�4��7�)��d��@�a=<*���d��$�
̬�8���N!�Y~�E�o\��!H���$/��!.�9���!F�V�,!��a�aדY��$�0��!��1քAc�do�[X�a8��9:�N�$��p&�a����l��($�!-w�!=<���4�/$�d�,�D�*�X��`��V��X�N�X�O�e�E�I�R�a=ėz�pFQ���Xm¾ߑm<D�a���C��}��7�;D��a��Y���"�'���!LjԪX2�ať�]F�z�,%���T�i��M��g��l�|7"�Ve���i��1�lM[���!���!L���43���ʨ@ �a�e�G4��U�lg�_P�a��U�t��U7�?N�E��m~]�F���ؤ!�,̪�<?d�n.I��!ť|���|�x���hP���բ�fo*�d0�_j"�$/�šRU�J'?߸�>-�-NߦU߯W"�|?W ��S����f��a��e����{�rm�B[�!�-�>&4!ױ ʪõW��,� �;'��e)�Hs�od%����T��,�A��E��a��k�=�����C@r/gɥ)��t��Xޘaͯ�1��''8��b*��|I�E�b��!�,����!�oy��Ԡ�B�H�P���b�h�A���,�!&!L�;�S��
"el��9`��^�}�x7�l�ĭ�'D@�!H.ݬX�!F�~�,%�VO� /�YFo���'Z�U`R�A`]5���uS�t�^�a~�r>��&��7J'&Ħ��0���� ���Eg!�,�!=�T��l����l��q��l��d��=�T!���)�R�.rz�k�b\[8�S�� [�:�!9�������m�`�w9��q��:)�X~!ߪ�8)� ��L�|շ�1�X�A@���:���U�T�T���i������gt����mi�����ՓT!�}�޸8)���Sޏ��!�,ͤ+!Q:�S�8�*�z%��d��`g��v�z�U��d��M��X�+��YX@�!��IA��?\͆R����(�t�14jx��խ���h��zk���lx��k���@�!��AA:Y�ި<\�:�S��,/\է�5���{��e���oP��r|]�ln;�ne�\�&�!5@�!T��9�nB��8�(��gi5��ɀL;�E�<FF������C�2�e���c���fL�.0�M��yaEo!��`1B!�������[�6��z���s�=��Pܗ
�=-M����Jv|	'������z��e��B��n(	;�ѩ�c�VW�ى>��@�0�'�[��Q�M�v�Vr��}�_�H��WB�-�W#�]Q��8��U,�!4��慜�a�f�arG�a���a�����I���a�c�!�,�!�$�!�,�!�4�1ℷ��X��&��T��m�mG��$#������pp5��aD(b��E�5�y���Pĳ!C����k����&�yx)� �T���O�����d
3��f��qUs��~�a���h�X 9ع�,��`�D��i/�	(�)}Y�֕��~��FZYN�n?j���,��_�\�M�����a7��l5b�|�\���>� #�/���:��ϼP�O��M�,ӵ+��R�C� ����ڏ�&����`Bd�6Q��q`�tB8F(L��D�+Th�h�P��GLzު{IY阘k�s�W��GH\ټ��(��Z[`Z�~��J0���Y��[PL"ε<y�ߝ���=i�r#'J��"M�$�A���6o�Yn�列�:��H��Y�LGJC�r�t�%fGя���5Ibj�L��V��8�'oc��\o��:�A6lT�����T0��Z���Q�[��.`��G����w��6}��2*vgi8rjnS�$�:���I�XZF��k������
^$��K��|��Ykk��7;�q·��
���zɘl��vh^% ~_l�%fC�P��=ڡA�W�%نOv�Si�<�z�>���*s}߃�d ��Y��[����w�>�\|}���3�"(�}Bb��A�@F'�لqk��E
*���3������.�6��!��d��[D�w�0!�ѕ��1�W dLu%�9��_A�7 ���{�ߏM�0���E�i��t��ji`:O��m?^���T�M�侪�n���/��[Crׇ��-l�7$�X��5��Շ�I��l�*�&@MŹ��)Μ�H���)w���7h���p}vg��� X��B��ާ�v��b�#�oM��萋߉���JL��s0�T�9k�"e@���č� ���<�D�t�U�kD;AW���顐��9C�c�����k�J��g"��d��sY�E���|�� G{�-32���N�0�1��S�!9Hi���6���g �&��uK*K�~ �9�\d�����<��b����h�.oi��4�5GЮ�O.�}���z�# �Z�� ��{!�u��l0F�֣�zُ�F�@]kO<Hp��ި�kK��2��>�%�I��-;\��Nx�H����̻-�#���e1�/�uR�ݟǩ�SO�`S�T��� jNi4��h@Qu{5��K�j1��"���1\�@k�����~?�����Ae��ßOS=,8�e�#�v�o<S k
E_	����AV7�ՇB�H|"�x�Du��ƀ��1��"�=��?�D��J˰��9����0&] �1�>���F��=0mY�n��}Y���0��=��_^��N|�b���W4�`�ܳI���yB2��6�Ϯ��w_#�҃�Mw���
Q��zBj�%��0=�e�� �jt���H��S�M{��B/t\���ԩ$K�S�����vm*��z�X�Ĳٸ}n׿r�ߦ��V/#�g�{��2��O�m��n�ن*	�����{�)�U��xE35�"�u��{���i�#_�NbjNo����_��IQ�`~��vn���m	����,�>Q��3���8�ـ�8�tHk@���-#x�݋b�^��ky��Zѯ_��}�E�KѕAǉ���i'�~ ��y*�,$p��6�☿R2�L	�A�X!�|&���qXT��\������]d����Z�������O�����i:P�ؼ)�=��|�U�.s#��V�}=?�#��s�	1/�����\��Ȍ�� �L9�w=�p7�?�mh1.;��^=D�ۥ�DC�'rqh���ڹ��F'�?&}�82!���	*���N��r��ߢ)}&���W�ˌ�~��/�a�ͺ!z|��\P&�Vd!����?�5�� �A�O���{i��_Aa��I��uj�GU����u�M�y+RP��7�aZl�!���-� }��
шn�ۡk"����bO��m={���6�n���i�}���	��LF��]�_��Ix�C/}��V��@�s�}sC^	�V�ha�T�Pƿ����<���=��/I?Y��W�-�YPrj��ڏ���bo{��I���{-ɲ��yR�hHSo���9�)(Z5��9�l����t��`������m)����'��	�#���Wn0';�]1M���b��<�͇?��\L�׉;[��F�^Ye��U2� ���7YV�d7/��R1@����ζ6�ٿ1��}<�,P��+M` vVEj�bWv������z�	�QL��c�x��gqTv��H�� ��Zә��������Z����_.\;]��	G�j��ZF�K��մJl_Bο.������#�����7>O�"��|t~[",DU�ҍ}pj
Y����*�Q���"O0�n(�A��G���S�t�֪��"����º�͓���:��35��=��
,2�Nc+�t�.�*�&�<��B<�������8�櫑0�����8����f���R�Ζ�J�F�Z埫��H�~�,����o!r*�5!J#0g�E�h��rY,�Fݽ���a[Tg�R����á�)�KX��ѳ��G�t[�� �#�-��@�i,Q��x�.ã��03��f��el���-��ڰ����o"� M|����
�`��d,湉xp�cj���!���|��`�����e�V!���s��e���NO�x�����2�"�d|ͽ�Z����>$X��V鰷�L�m�w���V�n2�)�T�[�2
��>~������N���g�[��%�?�'���Z��C+N@9��*=,[m���I��A_j��#2
*C���(nV�N�C�¥��Be6��=r���%ob�B�~�$�7l']��I_��Ҹ'���������3�����w
qP��	^�mX]���/���&h v�FTå�kW���;R?n+�ٶz&�Nlǽ^�B����
{����0���~j-D�N��.�r���?+x���Ѣ�B*H+T�>�1�u�^���A��˓����B9Az�Ł^a��tgOī��>Uֽ�mK�6F>p��"�Z�{��ƫ��%kn7��2׌��T�����?RL��i��l��/��s?�A�{�̍a�hS�*��[�1Rrl/�@u�֋�����ò�����"�x��c7^qL�F�vӻ��a]��r�-�tV͊m<�:)-�c-	 ������rB���+��I���O�^�}��ym���ή�5㒸3\�:��$Gw8%[⼍�))]�J���稬׀�L�����*CH�B=�j
��"�ok;�+��������b]E�+}��W��a}�&R�'=��އFE�gz��I2e&�#hW���?�/�}��sy����)=l��:�������AM��2��"�����:{�OT�7|�W�x�I*�F�`A!cE�N�O8�#?3��j���d���D�0T��u�f:d���)�E�gl�����+�
���!Ɵ�+�ʱf%�Mⷒ��C�xa BB��k����ˀhx��܁J/'0�J�H��gX��7�\�b�!�d�W�F�J�""�Y[ʝ�9�+!��) ��)�/d�6ވU���K;֨��܊��^���tK6�������ec�{;�?��A<��ׁ�A������()����X�ͽ��Ͻ	mU�Ch �?�i`�l���+$0iKR���ǝל;�=��U� ���z�&r�d�=<Y�w��w&@�Rb�8#ö�r"fil��6�_aĝ�+F6�swe�M�5�˭1A����~(��I5hv;4�lV�/c�O�˃]�Nj�������tڌ9U��VND�OW�Ԓ��F�y�^�d�>��Y[>�x��Ƀw�b� @BakU������I���ru׭$'�Gi6>���{��j��9�"`�WC����X���Jpݰ�%(2�OD��w�T}���e*1���TW��˟/������!�����e�Wi��+K�NQ���F1C6R�j-��m��%5��:�ꏤvpܾ�� #�0h�uȜ��Se�Ԁ����>ao
0O!�m�d�T�ws��&[Y�;w^
�9���Zϓ�=���+�6�\�����"R�Chچ��ߒ:�����Z����\�C�(1͵#�,v���|Ò8�5I�+�i j�/�߅1�G8�_f�>��kUBfw�j���ii
v�i�� (~I{�nOtqsx8�,�z<�a���Q2���^o����8�L�!�w�6�LV�G�.yQ0
���/4+[��|��2�s�Wb!L���q��k�;,# � �)�ŒttH`�v��n^�y��5�E�S�yF�(�U��^�������
o�-'~��U�vH?�{�&���8	���j�y��~l"�b�������ݣ�TӨ徫��%]K-��K��DlZj@����94�����Ysv�+>����ޫ`��&�� �+ɐ�Q�s�L=V�[)�*Y���F��ۉ�&\V'��ִ�E�^�R	{�桞��.��S�Sz��� ��}�64Z5#ա�����z����*�g�0x�<-��]�S`��v4^�4᧣.#���V��b�����?��r��2I���'!�ɞ/*����U�~������]�'�x��.������	�&r��,[jvN���J�h�WD�A�{ �Q�q���ʳ��d
N��w<��P���PS��(؎�-GI�7���ݺ(9��f#�I���􂡢o�ݱ:��0$�j���749|�,2�pj^xҿ��,�j��\#+���,<�qퟐE@��e{�Pj�!;G�W�y��}Cq!�?��m[���f�_0IX���a9� }����_��'l�K��,�!�$�!�,�!T2<#%'%#-/-#y*$#4R\c�jdcmomcegec�r|c�jdcmomcegec]_]#%'%#-/-#ksjpvmsob}f-V "%�("�A�������������������������������#lHcQHJdQU'%#tP~Q@FQFiJ[JFB%ks')+e�`nm�hfe�p~}ckfecmomce, ">.(JWBvSDAaLFL%#=w\OhFNFoJHS%'%k�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#�����������������������������������#%'%#-/-#%'%#=?=#%'%#-/-#%'%#]_]cegecmomcegec}}cegecmomcegec]_]#%'%#-/-#%'%#=?=#%'%#-/-#%'%#����������������