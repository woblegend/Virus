MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  L ;sI        �   �   �      N9          @                      �                                      � <    ` �F                                                                                                          .text   ��      �                    `.rdata  �F      &   �              @  @.data   �   P     �              @  �.rsrc       `  �   �              @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        s�ةyxr�~����U��%�1M�`��_�"�\�-7$ۭOk8�{`<��'(���n�U��{��dod>��q��nڒ�V������By�ER�t�b�|[�b�t��������޲#DL����}$�r!��e�j��<�ݏ����ޅ���m�9���oVEŗ���?W��	g���G�)�sc�G ��L�lJUH���9�.2p��+�E[�m����!_�R�o�M�����1�?�{Y��aޜ��^�y��^��b2���tK�Wg,t@03� �?g	(�0ZNGTwD|V1�`]C���fT��	���Z$+�m�r��>�P�Q���Q>qV�4���_Ya���.����'���=ǜM���L#���V�Pl������C`���e���Y���d��Y���]{�3���ݩ��~�o�������i��#�I,�6��1-�'��/�5�+����UK���b��1���)�{a�?����=��BkL�Ѝ�6��U�Ɂĸ	X~�����'&kImn�"
6�(e=��+E���tM[��f	��g�z�^Ei����k��"�^���� w�]��/Q�J��d�)�ì�s��M�
���q0��_�$R�&,V�N��WF�r��3Y��q�7�}�C��}�}�2�#e[��^��97;� �!s/��2f���
c��n��8�gY�1'w�J�(���aG��kK�[����_�-j�Ρ(W>H6.[2C���bQ���۪� 3�d�*U�r7�V�i��qW����̜���߉�A}��[*�C���5#ׂ��M�TՅ<�L�>��Kڙ�M�H����*P½�W�.��A�1q�m����I�Tz�������fD�����F��kڟ���[{�Z�l�r�
�ro� &�zW.L��>S>=:�g�űK��l>���"����Bh�r���=����ߔ{77�d�����P���	�M�ܒF���F�b�y�x#��/ij�ۡ����4O)t����|;�@K)����_�[�J�X!QT픹!��@%����|�6$�YE �	|Wԛ��g��_� ����]�m,��#�B���z��>?���L�;���w���*o�z�[g�]�i�����<c�}�k�Z��J�G)c�1զ�z��(eٚK��߯�C$[�&"(��.s�>l%I��:b�GiZॸ��a����h����U�\-�㒶9R�ǔ�c�j��nm�9���*[��P����:���h̬��S̜���k���~�5�@O����Z����S�	�� 88mmwL��A�P#CbT\<N�wS���/oͽMP��<�o(]�o�>�0�z��Ik}ʽ7��A�yb��oz�A��ְ�>�z+��&	ͶĞ��&�ϳ�r-��2�_��-!p�s���X�čm��C�B"�P6*/0w�q��&�!M�%1acT xq=[�Af����a�Z�F2x �8�D�Iev��|^����:LX�3���apNW�g�7�0�p*�C�St���u��%�rC��ϥ��|�8B�BZ]v^b���l�@�Y���u#4茓�m��鏰YT"nW�7���RQ��8�ax����
�����@�=��#�r���������K!O1ee}9w� %W�2w���F��&��P(a�v�֘����ư*Bjڞ��%�92�����u��Z��C����&��4�ɯ̒�Kr$m5 R;�[j������KZS����',���=,�g���L�>��̀�>��#��2��7a�x�?�HD��|�b���!aI/��>9����K��j�i��V̩l@uD�fϔ��
,��u*�s���6"��� � �oeQ�A��bӫ�[)9Ba��v��kǂC�%,��wxS���be��+Ĺj��������>�rV�5_�Lt[��HS_�-m�c^���DP2�_B*&�4A;G�iGR߭6w�B�r��@\���m�f}ܒ�NGS2��.Kb��`f�`���֘�&�䤄Cܱ���T](w�T]���i�pD�����ԟaowB�02�������{jw�y�rtC��\��˓����0@�����@Wֲ�����l5��?�����*���DśV�Imb��U���p�[��_�E�Q�rJo��:Cz|�gx!g���j?.�,��zJ��}2�5y@૔!~��Wf��?�o.� ����cWGH��(O�Е�έT���P=�p�����{7�[~�;yie��,l#18�</���f�����+'�3v��L��\�fbڂqߨ�F?������8�������]�U�1�nѪ�WK�:�.����֑���XО�2�e�C��<\KA�Vp�]��g��c�뺵� jO����̱w��y���3��~�ztm+�/�����"�z�8J ��x��1;k�̨@���Y����T���:[r�Ơ��o�;�{�F)�6�~#�w�nĎZx��M��4��dIt9�p��N�!�<�G�����tI)E�p;�W���䠤d/�M5]�f$W74�S��M�����)��w{����g?I	������_�C$���ْ��yG�`��j�;���h�3�
��Nj�"����8����:�$Ѣ�r� ��n9�	H��#�~�H�/=�&��;��1�ߵ�K&<Q��/wLP�u�Fw�j'�5�
�'N�;;9��v��%�~ν�~'�V��n	q�k4oS9�Q(�fW�>���,-ݡ��R�IC��h���`��>,7?ғ�x�����m�q�%�R���"R*<�uQW^���������WS�*0t���6���51��R��6� F�XuI�+�z���/� �ʟ��A�E��&ld�%s��0���B�8E�(����֐��i#e �1�R����UՐ;�+)�'����V��Li�T��y�݅����Ή�W�)�?����:�=����3H��y��}�:�SR�����2�k�m].�ǌ�q"se2����E,�mE��"�⃹��5$��y�Es��>�@�/�Ġ��
��.,h���G�=LGO��]��=]�aT��8��qy?���&���{���b���5#5psG�����G��� ��u��J�ϓ׬�6u���EU�����Q4���T��kʑ��4��Z.�:���>�/�'M��MMS*Fq��Ѝr_�<py	%�pX� 6��D+��N7I��4�|P2ʂ�
{)s��]fh�z֔l/��a�w�*�T�FPp1�~���a�Y���,�T��~�)8�A��W��Bγ��E��i{k���1_��0�(�����O���2Չn�@.�cv��������5`��ų�m4�N��;��4Z�CQ����j�O���Љڨ���6C��m��Cв���+� �K�6�0�x����^L������y�$���he#S��I9^�۝�Z@>�8������q~�H�L���	��rXkM�,X`�B�rn�u�=:���*l��e�E��U:-?�x%UT�Ҝ?�_Y��]2jێ��y6t��ٶCJi��Oʯ�7�p����h���8E�
�
u�p�טP;����O��䛠�����lMjAe~�H��*:!��`��N)�L��S�6�(4�(�_:���t͇�6=�Ko��ڎ��!���؜��.c�f���߬u[�*CXi�?�����^���Z&�b�9|�`e|�����ݧ�	c}�`��^d0c���^�%�ABe��E�;���O���&��J�I�V3��5�F$��01kj�U(#d�} ��}��C���a@������a���<b~?냉��EhB���ĉ��+:.��fU7�F�V���1�p4�P��řõ�,V��C��T{N̓�>�^�@�5<�0���y�=E�ėE��!�r(g��Y�6z�E������O���@-j)��w��w�����C�Px�p��G�pW��T���r�-P:T=>Ua��y���0��z<3U�ρ�KS�L��t��SN�h0;4�$�P��v�ɡ�N����Pt�A��u��,9}Ī�B���B��H��_d*�J��r	�̄�P���N��pI���jȶ+�d��NK���͐�1bPK㎝:��U���ݎ�E�:��v8t�"���M���>Ȗ(��"��JV7����Ő��j�t5���Y��b�<Q	0ׁ	�`h��akKǿ����>�T�Hj��Ih�����G�oի��zw6êo��)ܑ���y��ȼ١�姘�S8N���B�6o�4Sfq߱?�GfZn���#Йѧp�3���o�4�A�~��k91�G9�Qlu��/vc����<�{C�]��%�J#���7	��|=�ʱ���	u���i��ݗ[���Aw�����6�@�C�	���{��ki��9��S�т��s@����3\}=����d�3���}��Ȯ�m����-,�P�
+���6��N��%y�o��ﴚ(�#������Xj��m���h�/�\`/N�����2��"��y��
X����/��SD2�4eNH�r)����IfM�6�*LD(L!��8�teAf/,��s��<����ʘ�_u�lAC���װ�K~���GMK�����8���m����C���vHGm��b��]���P�z�Éė	t~i��l@8I=_�He����F�F:�U�x7�.��Q�G�7�ul�~E ���P#�S!����q}J�����k|�*6Ļiި�AX6�xib�T_Ec<s���`JR�
�4J�a�L_L0ϐ5B	��IS��79<kșht�����3�WK'�U$;7L�]����r1kO����Zv��h�4K}��,��g��T��;/�.ֹ�#��W�ݺ��� :Ɣ$�kP��卓���̍J�~7��	��;8=��H����ɽ���ڂcӛ�6�Sd�e����Z��EA��+�~#X�_��k�=��+ɒ�glb���U�7�@UR���P�:i��O$��6Ûg�Xܬ��~�����@�V��_��k!�ߓ��$� 9{�f�C�_�u�R%�E��0���Ao�@9��)�k@��;,�����vd�F�pX��>�c�Ղ�����l���y����Ω��Y��Ն�jF�L.����Ѷ��GG���\O̚����f�O�S̕h�)9G���z��+����(+��üI��^/���rdW_�0��J�;��e�G���4�y0�`�����1>�ߺ]V��(�el>o�J��02��(3L���5v��m���)P��o���RO���Պ��NA����e��L���ŗ�4m�h�/��垶@s/���*A���ҧ'V�.|K��m/�-DXVjH5�tǌ'��Y_;�x���n�G�>��^lj�ri^��n�d�*�9�{-�]俶>
��!y���h.��鱨���x���N�˝4�]���EFc�W��ã��ǒ0ھ;�k�d9� eo�Y]��}�y�Ik���"T]�0(��f�Q����F��w}����l�_K _U,��(��&��j��g5��+W�Tz�I&�d�`zn~t�ᙄ`m�An��V2���;�d�>���	5"?XeHPI/���3]��A�Z�0�UB�(5��|�g���Gާ��3���{M���#�D� �$D񏤈��c�b1�]]�xC*ch�k�x5���F,O��Ӷ䉽���\���D
o
��D�h���]�G1ԠbK�)&�Ζt!��&���J�]Z��'��L���io|�;g����$�E���P����[B��m����KE3�����;􄆵�L��X����" \��k���?�ͺHs����.&��(Z� I�"�q���i��x:�;�p���Hc�¨ΠE֑}p�=��U�M��Ĳ�*"^j����㳐;����(]`�ug�&
.B1/�ؙ5ޖ(��z�ݞebF����/{���,�������I�%FJ���i�򍅬�3�"o�
�3F�[��j_�� RkAv�h�]��jR��ge�e O�k*�ǚ��iCd5z�nT��x @���-ά|�r�J�V> 4�腹�ux(C5\�h��!������V��I��!��ʬJ�%�����N���W0�L��7Djqs$���6dV*V����XcP�nZ�5���*̬\l������o=��r����'���ݸO1[�\���V�R{�m�o�&(hbn����}���yHb�Вd�T-�- ;�o���u?��KI��Xi�!Z����_?���|Jp�ST^�7V��)���m��zc�vi0]���f����B&���޸`�������P��B8�"P%��'�c(5��=ͣ�Ѹ�*y%X/OV���0OFe1!��Ϟ~��G��зN	V��zr9:�r�`0�N��c�6CDc���jg�9�t�	��/�s� 
���[~�]M�V����V�l:WZ��8;��W��\$y\�HH~��0���wg�j�ߣG���C�tJ�����v�*g�L��<v�l��o�0�b$}�r�,V�#n� �l_~}�uO���)�u�B
v諸}X�<�j1�N<ęv�t�<��+\.Mq��y�o��f�����:*xY�+�B�IO������ /3�	��(����J��p֊^(�� YCΎ���q�f�0G��F�WQ'���K��'*jPd�g�����BQ˸���j�H8�\Bh/� �<y,�ʀ,X�7����X2銽��g	t�ymnm*Ⳝ�w���)Sw�I��YA8��rear���$e<}20I�(F�X����@#h� ٬^�Ɩ�T��F�x;?v�6�˽䏘&{v���f[�>�����}��u��)�uf)7.��XNF9�S#�<ܨ�u%��`���4+LEjkO��A���m�� ϩ�h�R��>k�4�Pb@܁����M�n�ayՀ�RS*(�2��a�{0%�':�yH{�`Xj�T6�N�S�0xʕ����@����j)�/~���as�+Mz���X����P�7�d�Ir�0�/c��Ɵ ���A�(��YeX�^B��k���l�#Ӷ��Ԅ ���4��l�>�'?��נ$"�����?!���q���`q%�s�B�'�˅�Ke�[�N��z��j��Uԯ�%=o�`��s%aW�=4~�z�����[g�[���x� �EH��ҁu�6������o�H�vvd^���4�Sd��G��.���;��Z1�d,Oք�h��W� j#�BVOQ�þz/i���q��GT�z+�.�}��@���!V����=� EՔ��
�K1-i�GV��s���Lys�0jRV�;O"��9Iϓ���z���d?bz��C��T���,�*�~F��4	��F!�l=�bI]��>���y�\ȒBV����'��m�^��C�4C\na&���-a'4q�b�A���Vg"�f2�z!�kX01G�6��2�;���27�>T�
�w�e�"z��|g�����w7�iewc��|�nw�<i���� 0&:3�.�x��[�AOW��1�`H�m�5�`��D&Gf�m��L-���Z	ή����KETn���^���K�p����ԫr�w�������!�Y���`� ι!z�Q'����D�����eL9�]< �9�,:҉�U��]�(�Z*]:;k�f{^�w������|N�$ɧ�:�V*/H�(����9��=�3K�.�Ӊ��\[�%H�������r�]/���������P%G]����(��0�Rˉ{"+��L�E?�!|m��kǪ�u����׊�@�gL��W�uT��sLhl[�g�Č˗�
5M�m�f��SR~ļ�_r�J�5�~ �5S$����:�q�1�&�%{�t����x��^���z;�����w����N��C%S��90�t�I���#2�T�A��Gؚ̀^�9�8�8>���]�����Jޗ�0������mqL<aa�]��G��|IPh�
�N����^(�a�� w��"�y[v�G�Ա���^W����*.K�d� N���"d� ��˺>t��=)f$��'�"k��O(��H�� ho�<�y���b�X�Z?O��U|�1�Kc��d�`��`��@�	H��J�����Ǆ�� N4֚*[�P(��2$��z6�s���
O����"{�!� ��s���=�N����"K��ux�;�G.7(w��-O���t�R�
*�������!��g*�\�BH�o�r��Wz�̞�{�����N٥�r�v^Z����hO	v����!�ФzE �+�_�Zc��|ڝn�c�Ѳ#}�g��~D���0�uR�h�M+�cg6�J�5��y�: �t1�N�q�xA�nc�NQ�rح&Ct��򈚇�it��Iʝq�)y�kb�{ɷ���=�b���>'�[���K�ۣ��75�-z�������(��5�?Z����D�\2���3��i�T��3\�M���{ɺ#Ǥ�%����CJ6�<*Gh/�T���n�`�Ț�0��-C�*�k���iP����ww�2Y����v�}"_##�rD����'xP,&8Q�=NH]-�֮���Ǉ��ݻ��J*}��#��g��u��x1��ߚB���g6(?ǯj�&�Q$��@���Ay+]a=v����bΖy�e�w?c?{�2/UuX��^���W"Y�$�P�a��Q�|��^�$�4�_D��!�~⏴�
8/!�V�3�x�l(F	h1x��_E)?���?�YF�� 2ζz@�Uo�����Q�!��\�����bΆ��r���ru�#H�H
_FQ5�a��²�Cq��'�V��ҩ��T����,��n�A����c���ⴢz`��^]���>�,���?���7����P#�@����A��8ZJ�T7C��>��K���`=��B����׆�Q5�@�</p�H��~���ܟMI�
��ρ�%E*q�J��[8�1E���Q��gV�yvr�+�p2��X<^������MU�Ţ&��]��4 ��"��/�IXX72.��an�:��OR�0I^�B|�.1��;0H�!�qW��6��{y��^����w�t�?6t�C�j7�
�0��] @eQ��0�iA�q!�#	�02�{u�I���K`~f.�6'cE��E�����K{��"J��_���]W�� ����F#��
��E�8��L�B'�fU�'��7��;z�*��M�j��l�H��z��4x�+5�u�8��֙��_\?~�cz��d-�/�����pE�jQ/V�>��s9�;���^�*x;�#Β|i�̎�s�8�䛬� Jn%�i���:��W���*55^�G-}f��es~���
F��4UVHs�M�o7Q����}�@C��M!f^��=ܼ���;�,
�	2|�T�7։�=�@�=��n�P�,�$~��(�I�~
m30gl�s�!-ct�!��	����e���4��NJ�i��Q�P�������A)IK�J�+sHƙ����Y�	�=G?˝j靷�[����Q�~�%�� �Q7ȉe�!��@�Փwˬf^�E�"Z4½Fú&�,>�]��sі�Y�ٚ�Q����o��󦁻<�:���A!�<d�vL�������*�
��ӑ||�����.}��{L��@-�V��OƸ<�{Ɖ6��bv� 
�ii�����ֹ�x�NЍM5�Ad��� ���a`�/��m̓�c�a2�+Q��0qf���Fkƹ������ޛ�����ސZ(_&�W�D5�lK�yV,磠��,�"��gX���ԞΆH���v��ם����aI�=@T,�˗#��h���3���!Ss�����?�����y��z*<w뒠i�0=�4��qz������,B��O�L��0vT�2չ�,�~f�í�����#������F�\���Aq�ކ��'T:Z��|f���8:�_���F�Ѕ���Tk�=�Ã���{����䰨"��~~z@G��O�iu����So ��|���n4���$LgSE	��WE��T	��{c婏�pc��������ٻ�`�|T��5�G�<I��{
�Ѧ��w��o�����0��<6�$YR�iw�����g%�+5��G��~�QG���ܼ�$���`�Q�����1P*Ѹ�!�h�ӆ��25³~��H��a����;@<�9+�l%MAQ����Z�9w���	o\��&e@���uC���.�X�Hh�����d   �dV4 �������P�[��A�0�   �I�	�u��@Hh ����4   ����P�[�����Ã��Aj j h����h=3 �j   �ʸb���O   V�U����E�    �E�    �E�    `��D���, �^B ��]��>O ��D>O �U�RSPV�U�a�� �VB ����Eg���U����E�    �U+U��JA`�!� ���+��RRRU���> UhD$ �   ]�E��U�a�d  �� U��EE�o ~��� �����}��ǭ�K�����l��
y��R���)B��Y�/��3ܽA���(���d����X߱G���Uā���c)�[դ���13Č��=��#��2l�j���fJI��������X�Q�w�ڢ4.
ë����Hu���h|Yo��_'#���F�F��3#̀���~6v�j��W���a.})b�Z�����#� �qo���@G0^��G\��>y�[fq�QrJ�	��ߨڥ�KC�&������TU6k�L�ýV邈���O9y��&�_�ۓY����8o��D2�����m9Ű`�;5��p"j���a��ծ[D�쒀���J[�g涾bcEEn��*�0�� �܁d��c��}$�Kj�a������3��g�q���_�yЮ������bN�j0��y�I�7=���cF�n���K(嘎FϜ����F� �F�X&�������qZ�ȑ1�;T��Mi�����,Ž_qZSEK�3�&#��n������y-V�{�$��nr0
�1�&���GJ�s���:|Z>a��J�<�2Bq��G���o�A��0��{�B��q͊{K
�D#π�>Z
S�y/><bA�c	�d�d7���f�JZ���'�<�"_��t�$SQ��ٮB��Q���޾�6x�>V��;���r��%�U���kѹݓҷ�JB��u�pe(s�!S�5�8jU3`���$*�iEB�����=
gy�f��E��|��%����'`Q ?Z��E�u �Jљ������ 7&�D��%+��'q����Vϫ�'��v�����,~qe1 ��j$�3L�Ѭw������ܔ۝�
������+hGdU��q]anh�8�vD�1���W�BG�m�Y�Ĥco�o��1�u̴��˔�h�I=�u�K�9�?�́�٨S� 
����Y�%l4�L���G��M�3�O�5��޻�nTl�7�{P�'t�-u/������,+	6Y%E�//�v���P���M��(��a��̾�2X�`-��l�=��ӝ��$-��G� ��4�]�C�^ь ��	I�6Th�{��J1�����f�3���r�%;��E��	4&�,cc�[�!��Z�N(�%�X��(���^%�^)��9��J�֮��r6�Xm-y�u��{u`0h���2��v��x�hZ����1���ה����X�&�n,����'3Fa��ٗtd�+K,z��ż��ʝ`F��O(RA��Y����?���Yc�?�������@�>e�,ʗ�骷tg�����c��(� �Vw� ��:0�o@�q��`.��WxU՛���c�!����6�ˊ�1/����3���vۺ��, C<Lg�أ@])�+��bxֿ)�!}���I��|��*ާ����AE�XT�F�]����D7��=)�uc��9D�}S��3��}8�.��^��|>�/�Z�<tQM�/n9��%��@F��Ե fb��!���=%`w�@o����q_���������W��}ƒײ���Kd)�;EK��;�r+��\_�kC�=y��O깟r��ӌi��Z��|�3��U���2lo���XL88(w��lL<����ٗ����d�e���Fۻ���R#Z��h�$�����H<a��)�s&����j��Hqc��N��o�>��B}�w���&�L�K�9.�D�A9R�M�K��Kc�os]�7ܗk[�.a�]f
}{����	q��t�89�̵�azv��>��4y��E��`��{���Y��N��.}�E���;�- �3��+�ݾ�����F�է=C��Ʃj��H��
ZQ?�7[����m�N���ۏ`�;��v��f�wf�Rxf���Q�`��͵�	�%���j��%���X�p2��=�3�����i��>����f3��L����'L��`� ȃ�3��s{�N�3i``�]� �O���WS���j�J�	p�k(Z�w�h�C��n�6��x�}5v���݂.HV/���]�FmF#�%5�_���H�����djg�]�G�y#���S��n�{�B��% E�E`���L���a21o���l�_������!d<X���<�VJ ��|RC������� FZ?�M�P	������]��7�G#󲒳/�|�`�u�(��z5����\

 \���7	��}/����¹J|~8���L�oůj~&����%ٺ�h��n����M�'���!���0J�&�������(�F�r�ʃ�6
,��P���HH�kA�0Q���f8�"у�j��]O��.+p�q���lc`	��~%2�1@��X�0��0ۛ��~Ɋ�U~x����JxR�q_�mxvd�	�x�H��-�_��qK�8bO�"H�w)�T����Z�r|��nǌi�W>�c�y�lg���ڋl�K�)��'�Ȭ�ї�o����|Y�dX@���m:�|�O'i��_�����:bsz��2Z���?[{0D���o��s���y�"��n+R�}��H
��L*���+SHY�M��"S��y��lm���L<�iR -�v8�u��K�'�N���g��[G�wߓ���r����wF��K�b�<��1E���(����|s��V�7����^�U��^n�C�LA*!j룏����\�Gq���b�Rsz�я�� }��u|R-�w����6� �-uz�D�a�ٕ�y��`�M?IVs�����������u����6r�N����0�ֿ%��P�f�nW��8uQ���[K<^��&gB��2���Tdo29�Q��ô�r����&�"�U��Ň�ߐJg��l\ 3��O�<k�ͨ�W���G�N����
Ђ�Bf�����}��Mr�6�1�%9� �1��}��>�R��~���*� 4�	}��L�U:����c���ʑ������,�2��*.gMJ�	�6��B��U�k�x �ͷo@g�O�P��0�9��dm@��5;��!1�W؛�g��愎�ŁW*|�Ӿ{�����4l޹�j�^�3��Z�7)��ʅw��%�g(]C�/Ch���y�<�K�jI����24�ѹ ��\��[��XFH�]|���L��Uw��	A��EMO�.����`�]((eM1Xs,:/���Gt��/}���������y[���Q�&��V*N,��  ��c	
��a��c�C�!|���# GXY\�o�JST��gm�|���@g���A��W�����:*�CƼh�3�QO�z1�l�R��֘�F�8HX��+�N7�ڕވo������l��X�4)�#?��~XD���ړ
��N�rm�ӝ�^���=�<|����TK_$�Σ\�bJ�,7��(���9v96Og��$����
�Sc}��̈́�
9CW��A&cw:5L~��xn�������t��k,��I��ck��~��{x]��O�!�	���-ZDרz��x�Fj�W��-���?�ЩM��A���3��+�$	.Y��iy���G�ȫ�]�����8�i ��Ur���\6n�D��I�:�� 
Nc�M5�@n��Y�lt	S��/��y;{J}\��3�A���a@='w;�wo��E|?�R�[ο��J�;�M>5�}"�/�ز��Z�4��̫�x���� ��p"2�\�x�� 86�54��B�j3�s�lD�,Ɯ�}�8��<����W���4oD�ҝ���T}�tn��IPm�p�.{^Sl�*���Y�P�S���h�	�J�%�< ����D�M�MJ�g g����x-���h��w*5�T���b⑛�����E�m��*�mH���x��������9�$�29k|���. �*8�`�(�#�֑^��K'�!�VdV�[�vB���@@D��q'�S��kH|��L����\=�k^c���:v��Gfy���W��m����`G��
|j��A:���@3���"�;����f>�e�`�Y^���/�	�������8�g���%8Rq�r��<���2��,7MJ��E����n+W�МI�����K��Gx\�?�Y{f��Uަ,���>%1�;��
)
b�#��=���.B��6>7L�m"�K'��6;B�L�����r�Ű1�#�ݣ4CJa���X��Ŧ�Ye
#ӴA0�k�6G4e��`f����Ȑ{~'V~yI� �n�#���1%!�,��<t�ηp��A)�W<�iԀ�-�M5����K�_�u �"&#�:����?��h�7����ɜ �I�w����ĸ1�A��X�,*햰ܥ��A,��M
��-�[��b��d�}�c؜��%݅��R�oJ��|���v*Fi����ar���g�S.�bpIR�3��>�%�lZ�}2��k$���{	��7�]�>�]�Z���`��	�4@��� �Z��x���cQ�>B��$����:�U/!ys��@������q-_j8�"H��Ϊ�����"��h4]�]W!&����CLҹW]���pO�W�l��h��B��D�*��p���#��a��P��C��F�b��r5����O>��jR�gQ����ڀ�0�~jRH�K�,
G�"+�i/���n�I�~c�~�
��)<*1�%��!��fr���b�?���'���Q���Bm���&�딁3��R�C��f���!��kX#���� ��K��J��M���&�������W��_v(��eZK]e ���Q'���*J���@
ȰN(��ﰧm�v�`[,�>M{�t��G�N��3��}��'��!s2
нٰ'\���������3W!6E�	[j��O�>Ç���"�2|�Fò��O?�s��%*pb�]@3��S`��Oɨ�;:N
w�c����E�2:>�O����W�ޟ��{���h����阒̊��6�em���Z�:���)�m��U��nzh��`�� �u�B��C�ڰ������O^�Y���jE=�F�9������[+��T���_kn�����r�޷)h27�)KxV�w�^���*�q�DE�Da�Td}�m�e�8��W�Yo�d����m������ ?pH$C^���v��������E>�w�qD+��R��5�4>j����D�'K��+4V �5Uxl6�[�w������Hϒ����9	�=�MPS�Cz��`O�3��eF �!��~����>�׺�)m�t�=9Ve����Ҽ��\������ӯ������2�F�j���˅E�x��ä�{{�n�U=N�n7X������o=c9�FZ�4�F�k�ǳ�x��Te+�� �L�Z���v���u�� ш�$p0�ԗ싞�����������N���A�xc������k���cE)�6����?��|K�(	����d�=u2�%r�H�
7��Fu��T�eSx�r�a�~(د<�`@��|�|:����|M��rI6�e��%�&���^�Q���G6��>{6����o�Mo�}3z����a}�h8,��)�.��Q�ZRE~1��K�=���H.���Ԥj����0�������}U�`#��� ��C��LEhg�B1`�X�#Node5dM��[����C�8���"�8KI�Rd�^��
J��{Ƹ���x
l�"�}L���C��aL�P���eF�~w�.ؑk j��ӊ��_[���n|����4AB�H�"f�G_1��J�c��auzh�w0)�����u��y����X��b�Uk���1�-:!��7/������ꗊ�*���~7q��j>y4�#DvM��%=u�t�۳����K��
��j �j-�`���%�z�)��jh���щ'ܢT��@#��JV(A�n5䢜"L�զ`�52�˥~��@o���v��%^\�Fv?{��W���h�Ƿ0>��z�m�ʐ���vq�k�T� �B��aށ.~��I�s��?�ʼx�p���0+�'���mbI,H�:k}hn*���'��e������Z.�SռM|�4��ƀ���� ���T�ʭŐ��z�)%�(Ht�����"
v��>r���8cF3Ê䃜|۫�z�e:)�5�I�+�7��S��l,����|yC��#���g�]'_Vo�.�9�h��mL�{���^�H?��I�~j+TC֢D�-��q�)X���dBy�Qdyc4���8Ձ��@�9��~��pϷi>Ub�J���r8E%Ux:�S{/���/�/�������)��@��@L�$~���lx[k�Jjt238�����x�D���T&�ZerV��2�Q���iD*�1�Ō_hl-*2�� ܰ��o!����*�9�;Hq�PX����AwɃ��Z׬�4]2�����',$�d8��+O�e�*�qCR�0�S>`��(�X4�Be�Nu�KI"���S��;�2�TO�Q�
�{�M]��p��aqF���4�g�<��F�P��p�+��s����M����j�@q%#"����?��sk-�[��f�����0��<�_c��JqFf܁(&�`huq��_7٣oz���'�����v�fs0� �d�v�"�,�]��S3{u�>z"��e0C���,ߢ���,�C��s��ܥ�F6���7�W���?��,��v��AoX�"ϩeS�v��$[yw�������^�U �$u�vK���3�Fk�gZ,t�U�n>Eu�P�΍s��R��'%R���#w������ �εlQ���^闍�|n�dK�Kf�`�1�?��w��@���-8dFǪ�@CO�I�b+HA��=��eU0B��c���}���T��X�F6;�g�s �-x"ʙB�n����тG92�^���?�Y[��ބѽ��(7V��O�.��޼mR�"׹a�?�De.k}�3�\��x����8G�%顤�>Y8m$����c����
�/`I��p~1݄#�gOB>�y�U]sc9_� ����y빆�K���"�&�%�WO������a~�$)��WU�z
yM�$�3�$���=��u>�!��@jh�Z7[�J#"L����t�"���<�y�m�:� azп�]�� �\�o�� n�6����M�t܋����F����)�9�"M����aoh��!ptj!��Pz�X�(S�K2�n:�w�wվ�w��N���YM��W-�~a��3%�O�z|�y;A��i��[[�^�k�L�_�ɧ�i��$��a���Y��]loL�����L��r2�dᕶ�J,�'��Ho���� �!���e�4����Oh$R�<�p�� �9�(qB���#�H\�s�v�iy+��fT�]�x̂�fħ�<��(�F���mD}�%�З"�jҤ	��fa���%�5wv�7����9`�}�l�	9�f^��h()�R�,�>K=m����E,�{�s�u��޼�]�b�`������[Ӂj>��
����F(A;�`����fQ��L��sC��a�ZA��jX�F�{������`c�аN@+�!5�񪯯1��G�3�����t��m�h�� #�۵�+z�M����4�r8����yAO��Wd��@14�D��_FP�q�>ӫzd�c@ �|1��T�5;ZDJ���H�ɺ8���Ի+��!e����m_���fa
�@�`r�΂>���N�6*��7�$�␌*3�e�I�@:�y���͡���� EX����U��R����<�I�'c��3O-�4���svy�s.��_л���a&�1�M����h�QS`rL��|�c�o�9,�`�lт�x�U�����V[eP�D$uA���ڜ*�a	lX�p�M�}��"ȿ��B�aS��3N��n{����H��#�~d�Ca�`D5*U�( ����'CLևL�j;��{�>��{�����,��D��39 �����vԪ��V�|1v�AdO/����3�Us�),������1Yt��Ӆ�:��gr�E�t�+������{�=�h�i����^�����.��O�B�G�~��?D����\�eB_χ��\�9 ���	~~��g�C���D�|6�
��;���=�Yu>����2�#��el?�������oC%��So1�6���E8�G�=����/�P����B]
r��C�t���?�i��⮯�D+��M�d�l[�w"�3�%�VY�
��&�B�-t�a1��+�-�����K���~��i~���+��v�����NWy	.t�/��OD=�Pq���{��@��8P�K�]r�2�_ ,�������P�<���g�(�lp��
�����9�I���D3/�����3��&�S��ϥ	��RSO诼̳

o=���M���\ۋ�3a���[�Q4^��i����_6A�1B�^<��;���E�A�4ܦ���a�\�[�˧��aY��0.ԥn�S� �\mC0�w�����xY,���������ӓ.��X�ݲ��{�������Z��@���~�i_��z qA�0��-E:q�J_�PQN̏k�r�-�@�s�w�$�l��ZJ��� ǝ�B@+��h�l�=;P|��og�z�eM/��߼�N�|I�&ﵵ�l0f����#�T� οE�s�'���}&�:���S��f25^Ѱ����Gunj6�H.�v\"�6�?ܷ�Q�Ӎ�՞�FHw��Nm�����&nOG,n)hـ��q2(	�랢.�ݻ���d� ��7;��a.V�o�(k�'%�r4ヷ��`̙�@ɖ[� o�Ș�\�-\udE��+Nn��^��n����&����#��1{�@��~1�~s���9�ۖ�w�1r�/+r�Ϸ��ҁj�B�פ�[�Q��,�K���.6������V�cn},V�פql��Z��HQ%&sYb������ IQ���R��*Z�me���|ᡓ�e}�ʶ�eCe�m����t#�%�<�a28b�t�r�����{#����ug8T���@B��S��k'����)�}�J)8Y�S'z#(���J�֧�;	��(��u�
b+��L���	<)C��)˒e�䰉*�Ӕ"�w�C���\҂�5
̛~i]v��e���q*�{ٙ���K�E���{:|PP��+��T<i*��$��l��}b}p���F�{R!���@��*z�d�A���lé�#�MEhbU����ϟ�j\C[@�m�W��[g�Dɇ[���7T���;�2����~r���;c����w3��*o[!����D]�,�a�"ӣc:���
��W�ax�00��'t���
�V��x�b�]���[�U!g);�'�a�vъ�g�8���A�kx�I��d�;�<�0�;����.�{=ι�=�����i��&Opҩ�[`���1<pzd	>M��?�wI���浯�	��T;�h��dź�=ө��W&=��Υ���wl���E�f�F%����B�ܱ�awZS�RpyZ�����u
���e�}R#�/����1�.hc>MHǗ�s�pX펱Zv/!.�|��}r�z��'j���� 0mv.����]YO�����=���������Bɣj�ްd�F�ǰF����&�sJ�֜���)���Z��ʿ�~�&槮G-"
��V7lљ�����iɯ0F���P��x���W4��F�~m���YFQ�A��W�k�f��ω��Lߋ��8 r��� ӝ�(c{T��/�V�g̾8��5P~� ����T�Q|�[���Ŕ�<��g�"b������q�
C����\����
G d���ְK�+��	ڧe/TJ�h�IX:p�v�d�Z�Łqؠ:������n�jը���چ@�АJˤҘ�u�(t�����oޖ����!Sk����Fq'��j�� )Tx��:`_O�j��GD���F��B�,��ufi��d4X�؏0.�X��,�J7�Yʭ��Mw�����!���@�������K�I"b�R���J1m�+Z`~�|!Ծ3�M���]�j�Q��[e*���D���(�95T/	�_u���@ӘN�o�@�b(Ҕ������&.�R���u?���� m���>��6��&���z+������	��Pe��'q�H*��"�����0�HNi��=�4��Z��?/���Cs�WPe�S�/��������y�nn";�F�i�:�ۜ*|��WG�Bގ|�<����eE�D��*!�zM��=MK��ܻ��i>��e���DGP����ţ��������z)���ɛk��Z�+�R��23;��g�J��ߪ�a0(��z�;H��#&�S��2.�lY�d���V����_�E�b=ߴ�EB�[xɹ�~D�0.+/V4�g���<s����z�qg^W�^{�:"�	w�,��0��`i��$�����w�;Մdr=����b8��0�A��Zf^�5��g[8����}�8��ﯧj��F�u$���ϩ�����o}@�(�|�'�[�	�Pv#R}�L�'�����
�wܺ�wL��y��'�$.BS�:��|�B�~7�̎�q�d�Vˤ[����1f=2��T�e*4�S�-2 �iF�jw��	�JTA��lB��E�G�LMܻ<�!L.��Ňt� ��Ke*�QbJ`�(,<{�hu�A�C����^�vU��9�>cSh:�i�J�+LJ�p~��j�g�<*>�]d�Ҵ"NZq���"�l���QE����[bfӾ4�/3��m^��g?��_:y&2y��F�oQ�	����Tc�lzV��*�d P�t+�!���V�5)nQ/$��ɘÀAoT�=�_`�v�-l��j�0����,���R�E]`i�s�#�b��$3��sMD}x��j���>)e@3ʚX�Ԛ����|�QZ�ŌW�j+&sk&@�_��u	z����U�8	u"^��6dZ������iX\1e5�ᄴPú�i��/�$^��r��4%��!���:M���PGݓ����E`l��xH]w�ڄ,�8��
�Vp2�uF �D;?DC�٠�j�#�[���hW�Vwz���H1U'������Q
��-$u��r�!���J��d��~�D�E�ޫ5���D53����A)�+���fLݹ;c�YY@�7�Q�t	k{G<$o�[{��SZ �;W�����N��+H+�m�!�`�~��e�0�PD��R�	îqX� D�4�Ad"8�xd���=��R�G,H�`�"#�����G� ��Cn�$����{��6��3�|WT�hg�M9}fGG
\��nilփ�Z�6����t�le��F����r���ZO�o"�F��+�D��ӱy��o����R	n�ԝ�q��~R#��@�2 �#���l���1���!9c1d.ku���~�88;�t%�`\��l���,��Hͷ^f��Pn�k���I��<�6N6��"Q^3o6�0����6��d�>U���#Xw�����i�]f�/�d.~N7���.�C��6�"�m����صJt��h�r,g�n����p�p���we��d�ͧ=��`[�p
s�i�s6�I�D��Fʬ� \'�6����K�V0V\8�I�����-��~��J2.�KSP����%Q��2�7�O�y��{�m��_�޵�U}U>�XRF�̷��Z�A�Tj� ��2�9�٘��"�#V����â���u�B�= �c��?����2�`y�154;��#���'f�w-\�-g���jY���Dz���D�@9�V�{�r�s=�W.W���kk�C�{�<�ƿ#�� �k~����Q��I_p��Sxޫ`�坁	��2a�`9�)�s�(�\0�y��q~�3/��q�$�ۍ����'�ɬ��R�;�+��|�����"�����P����۠�f���8��D~�0��~�~ ΄ʤJU������LT���dL��E�����/C���Љ!O!#��S�ж"����	R�Q�R��-Q`6�6&�f*r�U^J@C0����K%Y�q����5��f�fsq(�w��Ϡ㖊6{
���ݼ��^�°3#��d������F�gu�m������:]�dV�(�

��\E6dN��:��a��N��~+,$dC��Z��%��1��e�$�DV�L�-��z��Io'�C���?"��!Ͼ(���\��XL�ao��yu����mKU�1RO3�"��E�ɐ���@�]�wk�^+e5�^���^x��fX{��A��'<������h�m�MìJ)I*�s����C���_ܙ��ۼ}���3�wB�Rk�}EF1��ݡ�~�k�8���e��P�9�
V�����l�0�(��)�i��gْ�l�Υ��j�.\d��̻v?WkR���)��}F�G<7�1S��i��FG��ʛ��e�U�l��#�3�b�e<H�m����|��r�����l�Gσb��m#��8tlv�j�U�q�w���q�~��5g	%ݨ������0�������Vם
��}M���8)l��ZьX��fۉY��{|�w=��t�C�������8/��L�,��A�ŉ��	N���I�	��/���������d'&ϣ������ݦ��지�>:2?���f-�R�`:�=7~�<ى��'~#����2��Z4oByjFkK��w��>�Za���/�T"x��ϯt�oۤ���W�=|X����ɟ�*���t���w��cj��e�;Ҍ�Y�L]��� z����%z{خ���
��~�Ɓ�CxF�@\:���R�d�O)�Z�[�茒����uC?)"eg�ViK�{�`?�b�8���B��u�+�^�X�W
��t�����m�j�b�����4mY3��`���4��:(��WP��w�f'(f�J��0
L���oa�V�0���������zΗn��K&��R���B�Y��zc�����19)z����MLwLk�yS�ɱ��#��-k$kM}���1��6b(>�ϣ��'{c
��x{.��B�!�N����n9H�bW����c�]Yd���;Y�Wq�䕝U�CӁpe2i���e�[c�9�:6��0��|T+�?�˞��g"��C'4:���T�r�"�Ad\�Y�:6�	�,vߴ��u]�ș���ǻ���P�IO��K��J�Z�T������l�Ua�Gmv W:V���3�נ<�$��ʏ�>���rl(����<�.��,Ŗ �9L�U�,6��]��*(Sf�(�ޯ��3�qC!N)��z�t�Ğ��?"�}�.&��y�t�"I�p���|#/[�4�O�&��P:O��I�Rчsi?Rx�#_,QY�~�n�?fmpP���6ƛ"[̶Z8�mۘa4� �m.l:�.�r��Ѧ�}�5������e׆B?�9��Jx�5b�H䖤_e���cAz��u��P�Dc���/�lK���Y�eWaKd�����a���v��+-����Z΄.�9 A8-�+�2�,;��&qbE�@��ұ"�;��!0�����@���4�('��%v7-\`jxLJ
n��f�.b�A�����i�+�gd�T^4;�OC�a��sO�zR�܈06�����S>o�>�f�w���$X�#E?H衞i� �gӱ�ʒ��(�������3@=&���C"T� �}�/EV�2xEK�ȉ�DT����k	�ܝ���w9K�N�ݹ5��~�	�x���I%���
Nd�1��|Q�O7S���j�7�S���ç�j�c!�#���Z[�̫_��g�*���ɵ��L�	����0{MoW̩���5$F�;S�/g}]</�e��-�֟�z�e��j��qgT��ېv˧`�ӭ�����tKC�i�p�.��"W�^���5��WY\Wy�uڑ�J��h?q�*�����1"U�,a��c�AY�F���7�|� G��d�E�����P�z3�9�!l�J������N���~��nq����]8&���򆼼h���P�%%������QW!e]ʦ�>��iZ�r��� =5�IO_G�i����]߄:G�#:�;k�OW���V�[y!d��`��Z�[7ٞ�".]9M9~�v�!6�*�:�5���5΋�}s�*��4��0M���y����.AT��PoSȿ���@K3 ��Ą#�ת-=s(_��xZ4%OI<�7�7՘��`�H�e�G>��j�8���w9�[��+��r���vkw�,��L�ь^����,��pռ�u�C���/��w���z7|�!�\%O��v��l<#��ů�F�g���D��Z-��M��7�(���>;��4�Q���\XY5�V��d�N|�k65vC{ܖ^ˡ�V?�>����#_^�2ی���c	e�W��Ku�_ٜ��͜*Gc���m��Po�Rxix�0���!�r�䝶e$��K[NnUض8�ƅB���>����r�-� �0�xa��ۥ3Oa�"-�C�v�A��׈KT�}��L���{>��3ô_����%׀��0io����Ύ;g�+��K\ 5u���Y!&��>R}gb��Ƀ�A�(Jo����(m��e��:&F"�5�,�� ]����s?-�-B٭�&V~�|>���y	r�7Pb��\�O�e?�j�G��9="k�����*Z27t��+n:١e��{���V���	�K�";���u	s8��ll�\� Z��q���%]�)7@fp0d�����"c���,�I�%�ek91"c{X�=�~t�^��N�ߍ�K��q� "�i0�ɋ�Se�{�)f�#�[E�7�t���;�?͐,��\��uQ~������!l�5�9�Ņ��y��g����fS�4!O�:)����Mqϭ8�ФD}�;t,��&.g!�&����+�Q��o���WwlUl�&/��4��`	((Nt�(��@+��%W����?)���F�V����K�9/�@�8
O�g��i��F��Iށ�r���~P������zڝPkě�~�� ���BjI�>{�4�AW�'�UJ!�94�A
��NU���m���4r�6���ܿ�d�x����=��E����>"!�z��I�5�\�����'��#�Fv/��Ly�����x(�o������t4 ���~�P����������-3�7q�a"�i�4}Q<�}i�h���P-��%�2Z'�d�&B(�6����T�2��	������2�M��E�1p����u�������[��"�	���ᤂ-Z�~�p�Jm�����=���;��4�������6\�&�@���^{�qЅ�$����~��-^��ڰ�+W �Og���wk๬Eo����D��G¥�=��wn�V�Rs!�
���Wx��r����V�R�)���KH�+��-VQ�~xv�~q�vt�˻�x����tw������ΐ�.u�Xo���o�&���R����B�����Bq�((���]a!�G1q���6@�=hw~�*����X�KlV��/��L��~�_���/Q�{XO祕�ne۸C���zg�@�W0t~�2�=�On����o@:T��X�\��� ����Qs?�����>y�l�u3�4�nʫa�@iir)�O�u�Nj�HH�u&�1̰	W�,���-�&����-$�Xԫ����ߎ�~;>g�
�Q�=&�������r� ?��JQzH������j��%l�k�r�q�ɦ'��^HNN����� ���CL75+��ǧ���OC�(���i��`� �/��z��ˀ��Eϛ�9��l-��]�!�
��-~���h�����x ��(u��kIi��]����bWS^2��v��a_�����	�c��z��Ƶ�6N4��{}WQ��$��hW6�Ɵ� ��k�O�O�9���d�'�k��G�]/�_1�i�ѕ�U��K�8�=��pc\un��vڄ��[<2�іG?u�H���"�iWTE������(�~�#B�gzP���|�ylE.O�~�w���l)�r��s#��"�T�����h�
�Z7���~	�%0�#��!2�Db�T�Y�N�',ӡ6ܨ���{k�x�L|��N�򢞫)�Mʋ�ѷ� ��X�׼��C�3�D�����8�2 �b�Xū��ŉ;
9m4:�7�Cq�q�چ%}v�z(~�X.�"ׄ�Ā�/����e��b�����j��\��ޛŗ�m@h�z*n�#�#B�?D�뾂��h�c�ct"%�^�xr<�,���+��HOOѲc۞���3�m3R��N1 �q5)�]_��=+R�u̘z��\BM���H�AS����Ċ�悡 ���J
��B��*����r�vE�#@��b�Zc&N��Y|�����o��٨��e#F���n<8+��lU3me(
G�-e���JL}]�{�RR���G�HV��Q�'�^V�hfԭ��$u���PY�Z�X?U�b\ťs;K�+�"�ڙ}�½R.�<vi)�,li�rQ���I'��a��*��g�A�r��	��D��u��I-c��ٴ�X��)��f2�Hގp_��!��X���&w��t��U:���)Әaց�����YM�&����?��<�3�����̓§����̺��� v�E�s�
��I��e��*:;Q���R9*V(�R���f�=8I�zUO�p�z�Ъ���.�]��x���jj�]3�z��AVs!�6�����p�����ŏ&�.�N�@�	�
o�ŀ1�@_�l-����n�n���o��~�"j�
`ݕ�BɉxzV:����u{kX3���@�U���&H��]R^Ѳ���ɉ�W���+הW�ut�f�z`���9�=Ɣ�K��*����0b�ƙ�8ib���*�a�OR��8�l��3
m{�U�e��`ُ��Tv�p��w9e<2�$_J��I�'�2%���:�s��h�xY���`�&�Oq��T{@���Y�[�P�2>���@ D�P�wo)B��~���妊�v�?=ÿ��)�<5rg����fs�{�����G=��u���Y�3����Awܐ����ޗ�Z+ml�gxY��?Kf,�[�Q[�6#WJL��"!�% (���w����(��[^.lx�925$�
�xdb̛]���1bҩ,U�;#￟,5`�bNX�'w��\�H5l�mcۏ��U��S
��`��e�fYp0{0��$7������N�%���a�m���	����5�Y����BM��F$l�U�$<�f1��ۥh�w�0�p��+�xԿN�f�U��$�R�zr@��bA�?-9LĖ�X��Q�C�"�g���Վw|0D�&��<�o<�V�T�f�|���է�<�E�B��[�D��&*�Йn��vɳ�}T��3y�=�V�����A�����N���1�C��@ ��i���r��0}O"U����8۽!"�޾-4�*?p� ? ��RU������B5��߻�Y�/-�m��L��2B�y�Qv٠����|���MщɢʘnI���,��¯�Oq�eJ ��,�u�d�'mq2�e���y��>����s�����08.���8-w�X��~'�-;M��`S(B4h�#vVc��'v�8��dT :���{6��(���XP��`��l�V�Z���ir�L����04RR֗�x*�ie>�,Ui\LB�5�檑�L+��m?@��C�;����E�<N�(�y�Giz�ܰ�I��%���4�?�\��D��Z8��������'ɽ��yo��hl`�=�����ǣ���Gg	c����'Vis�s��(�ВB·g�F��X�­3���ٵ��8�q�r]��t�.��xM�K`�W#���_-TǮ[��LP��^g�	�8E�?R����?�"�V���[!R]�J��Cd{��!e=㥙^�
���ׅZxZ�	�^`ϛ>RI�:�;{��m�J��TX�w �`��zr4O��v�񕻚���P~��p|�}9��{�$O�xZz��}�7[q��n@��[r:�� ����g�紜��r�=�R�I�A� �ɧ���&@�[�G�AvB���Ţ��.�g'��7�fG+�^��� 6�u��9�?�����L\d����-鏙0/����~�
(NC��h^��QO�9ď���{A|3�U�J!q6���o�p�Bv���C�i[�$���F�0�4��OM�������Oʾ�ǀ������(�"���j\ϥV����L����1���/S$��R���Ϸ��c����e�U!�$�Hg���;8����YO�z�M,[t有7@��j���]��:&��d��<��(͟�&,�m�Ji����ˌ����ȩ��F+>yB�y���<�yf6O]'f�2�H�K���TV��.nI����w�^u�"�y��K׊�����NڽD�l��Yb��dv�א�	8����ߠ��)Sd��^������7b�	Hߧ�oQ)j�'��^O���0�N�w�u�v^I�"+" �F�XG��77�����)5+�;�3��#2W�@��D���-��ߝ���=luںݎ>�z�b��2_6U��^�W��q��Ro�r�u�7�K�c}����d�,��蛮-��n��ܱ�L]e���c��4�?<p�Z�u����t��r���-"�`W%�@����������V.���p�%�Xq����ҌN����E�M�z�����<��p�8+�@�*��d��|&�9���&�&�T��=�V-W!jT?ķ��p��'d��a7���	G`\��6��Ag�1�U`�<�t:��	=�<�VW	�]�[>?�x�3��f��ϫ*��OƳM٧��c8�J������̘�Gj^�7��!���:�liO�u�҄p{�X�F"-.�OT�_8�:M%�絭v�g=��Ğ�ۘ�]^"�im�v����x��=�Y���ݱ�����&��,��vC'o@;�䦑f �Nv������M�- �{KLs�Xx��B5�U���ހILl����¥_�AV��
��]'�q$��� ��Y�I��짎��V+�=�Y�۴�L�=m�E��ӪG��>a��*�i�|݁�B����J�r1��z�Z�K���R���7C�-�N���{ 7���pmZ�h��pϚ��<�M����:Rz�m:����9�x$�ܕC��5����cН���ˆ���$k���%�\�yW�0,��-�8v��J+ОjT�\swW:�����G�b�?A32�J�}��M8^�{�#���9��$��I*|�ۓ����^����%�Z�B��ö'�a�6���ˠ���Q7�~���l;��iϫ�6VE�Vע'[����e��q�u��M҈$�m0	�2!G`w�g$����]pjX�Iv�݋{̼��#�@2�b�.,���������rf�}���Lmf	�D}?�_Y���{\�㜰��~�dA�~VBHz(>"�xRUcQ`w,ذ�5���a�@�YdF������L5Rp�QW�K�߽3�H
��U�֔sY�b;�H��`_.U&9S�<�j�:��0�B2�%�2ɚGg�iDOSw���6��Y�$���:��O��zXGvs걔���t��[ym �r�g�\�Ϥ]�π,�)�[��1���J���:��Ē/����9=l�*�,Qt����9ئbD���P*Gg�uz� S�eKb�x�K7��w�Hf��fto4��a��e�l��=a�T�1]	�W{�"�UPK8tZO����.�fO�@B8�U��g�ų��Nz[�I'���AN��u�V�|�4*���^js ��U{Aد���,�Ӥʤ�V�����v�>U��ͯT��l�l�S�7Ɔ����t�W�0~FE�*}ͥ3��犇�����e"�F�^�G��߇+��o�c���we��N���<I k�M%ɷҤ�:�_���T�t��u�rC�bgIwD��y�Z�W�.�Z:u�eߋ�/�e	��I��H|0b���d8y屐��3#��u:�nc���+zVB�?Č���9RhR��>6�w��\��x�0B��\�L����is���Z�����b��+ǰ�`��.(C�/�Wm�#`_XM5��6X�>?b�tI3�U��I�s�V� Jo_=��M0�6/:*�s�� �S��(���K8��>��8����Ew/ێw<�FQ�K���2�VcM��Lh;8�z�o	�+��{�r[. U{��R�rΏ/�*3�6��OX��S�w�L�+n�Kf���]�����<�x�/�7>DGF��15�����,6������i�?���ߴUb.��sx��7*��
����&��UP�M[=�9he�5Ak������:���$��N%f�G��N���TD��ek�x;����}%�?e�<�R������h٨��N�22�ep�:�u�\u��@[J��(ȻI	Yh<��V0b�L�5Q֖|V�}q�7\��q/���j	�n��� <��O8��+�/��(ؐ@	Ke��H]��v��I=0�����Itv�0(zl��hUN��v���B��p��9�
W"�7ك�����ƽ��q�<�f8�#�*�����4����X'�����̶8���A�s����xl!�fT� .���O4��"�e�<&d^�4�9q<��զ^C��,~�_��H�D~�^���U���y�uVj�5iUy���o��b�`L'�pL�J�A}ͧɒ�U����W�E�/G��А�>�%�&���?���y��~)��?�z�rk$�fN�=r�8��mF
VL��?��hA�y�p.Z }��K�b�7@K�����#�3���,�L�u����1�<;"#���������$�~���'�V���Eۼ�~�:إ�}`�u��ș�"I��c,�cvV�	�r��?kץ�7[�p�.�%���O�
��J�y�b�N�����|�r����?l�Uo��恬Y�ӯKKJ����2սY�Wol��~5�b8��'�L�_�i���M����kx�� $��g��s4�Y���+��g:{��mPo�fn��!ۙ��wr*��t�,����+KL�j�� lg�e���YKQh�G7B��d�X)���>A� b�t|��	�2�Ģ���M:N����')�d��E���H�zԽ���kڟ�R�x6VKZ�¡��u =o��%%f߾��B�0�8,���^��(a#Խ�ᨪY(�p�sE�L��E���E�����P����86:6�,���(S$���6Ao8�Jǳ�n�	Ƃ�6�{&'�0���.����M�đ�t:��� 3��NЎ�(�XFR��`]~�w=����E��Ұ8���[+�.��Vr7B[�i�fh�y���>Dz��9��=��Ӊɫ�%c���Z���h]�9P˿л���D�f�<�qٝ_m�C�'iYؕ��"�3�zۋ�_��9з0�ݫ��:;����y��Ul&�]}��V���oA�/�/�� U��~Xv���㙋Y�QѠ'ߝ0�~,{˔���N��M����7S�|�����
g'�+'�ńc�6����'�G�F�?؅u&��,`}C����	���	;+<�D�Xj�_Gn��OI��� (Hձ�3̇�H�-����6S���$Ip&�(Ɛ��A}f��2�-�,��.'_������YT'AԪ"�vAG,2�m�#C���h�����$���Q
��Ӳ����0�B�h�'�l�wd�

>]B5L���
#���p,���J�P���(s�Gt�UKW�v�v�R�����!�`ְ�1y���ޕȅ�NC16�la��kkl�	29�Ѭ����9�q#K��n��&?�ѺZG
������'�y�k��
�ѩ̿�^��5���v�/�g�0<�)<g���/3R
Z��hm���ɯR�ܨ3��Cw����z�耙~dx�Y�'}\�t�E��h�;����}�g�ǥ��eɲ�T�RC!�G���$�i�b�͓���B����A?�jY������|����-�ߐ�+J��k�������?�h��Ȫ��S����yӍ�����Ϝ�F&��<��$%pF�aaVX}�6�o�\da.���V9��@1f��O�!�biz�Q��=Q�v �؟�|�����Ә�l�����`�Lwz�=��sy���T7E�@�J��4�Z<z�6xj��@^�"j:��ϦU���C�)����i9;�Ջ�#%>�,��y���Q����C(�� z��2�V�������"	������y0�ll�bQ�`���R��y����99�m,��;5��Yv�ЊA,�4
μ0�^V��bMVz� ����S��xaJH]9|Aa_�X2�LR\HԤ�&2źy�[�?q�ej��j�A{�3Nh1=��4�*$�х,�wc�,A-�^eBYxAyd����K��MF�̣�w4��I1��U?����ǝ'Tc��f�1�.ڙ$ж䁌��J��{g����>�Y�[
��^�P%4�ٚ"���g\�Nc����y�����۸�^�=Q+	�;=��s������r@�`��f�����5����3�a�u����+dK���./�@����*$��E�u�J�w@Y�z��v�˛bU�OR%��Y��2�!I�Ԙ�4~Os���`%W?"��T�H�&���?���F�5�C�=���|')a��z�VE@����iT�m��C���JDk3��\j�w��YY}�1o�^v��q�^ݛ夑��e1|�u7���zu}�r��9U���ե�B�@�3Ub��[�l�NևLD48՜����x<�H���8cLu�%w�T�P����ojsn������m+ds8���o�^l�^Pz����Y�)��S�ԗ :&K3����vz?6�t(^��f9!>�\d�0�D��kG�6�<cF����1�D9�a��ԝ
C1��ʟs�`a�����b_7\����&$��;z��e���q,�$λ7�@��㆛�����lk�N�h���\~>&���x���S�c��HO}��[h�L�K'q:0D-��jTPE�X�rO� ���<���@@��9�6{��(/�R��f���wi73��T|��ru���P�G��K�%�R�f�n�&3�*�)�@���_ ��������+k���c�Aj��Y�Ic��b��M��l���&g�Z��A�8O�g�O;ST�^�������9tV�Q�i]�Μ��(����K�ߋ~�F"2@6yb��Q�:�ɍ�g���|&��	M,��qe˅b'�﷍{3����;���m�$�r?D��_�����Eo�O��Н}lU�E����fC�x'SH+!���J٪Hw��e��*�k�P=��=��R`n�����֍0.��_���͖�m`�qҨ�b��$�E��[�C�h8��8ކ݆	؟fk�d]�4��6�t�[��h��#�����<x@�~&��q�y�f6!h�H?����g$���r��8��#�e���.*�ァ������΃�P���x}']�[I`2žȐ�X�ʬ��{�*�Ȳ�z���]G ��`��k�sЙ@I�umrN�?�4�D�R|�������D^c͇��".IT����o
�e��������������Y��&�i���Hxb]�Ds�C�0�q�H%dlN ��i�*34�X�=��`���V�D���	��ʖ����s��K� ���JY��.�7IM8�]��2_�;�PY�fj�o�r�%�Qe�«�oǅ<��Y���le��K�;�����k��S�P'L^��G�O/��J�6=[Ub���d!4��o��@Ϲۖ2O�������C����c}P6�2��vg��y��!�I�w#��L��1u&���֣<��R#�-f�4!���M1G�p�R���2
���Qd߱&Ì�D�Gԓ;(�㽑'�L�7�k�D� ����x; ����?b��JF�f�N;��ډ,���oUow^����_$@� ^��
���iG;x;^9��efj�zJ������(�o��6d ���S�?��U���Z��9e�{�A�O�$�לE�͸9�̾{Au�������!����� ���ۡ��l��e����) ���]���c˾���4٭�'�E]���/z�TC-������	�y��0���C!R3�Pq����(xJ�[{*$9��F��.���q
+���$�4��"�(pk6��+4��)�a��,���M�*-�����i0AX�W
I;�y7�1�ˍ�m�iGי�xÁ�F���p��+�S���3sl���b��)�=˰��~xj���������I ���ݦÝ���`���#��{�����.����P�N�r��S�� 3�[�^x�!��t�hb���e X�W��`,N�W�Zd.�.f��^��Y��h��� |�r�ÿ�B��C~�rh��&C�L�+�i̤)�>�σXoW}#,=W�J*ޯ9�3Tq��X�
5/�'�9�el�q�b���9��Ձ`�ʝSSM�P����L~J9�����.K�6��ȊZ����-��ɡtġ��jF�IQIS�C�7�<�?Ƭt �R�9�v���l������ ��
��g���5�>��YG5��By���ٴqhT#[��ݷ���,!�3�j�rM�)� \~M��e�60�.C��syr�s�b�J�5�29��#��H���� ��Չ�:������^`6�l%�9���j�R�o�>1�Vߟ�8)�9=�`�P RJ�1�4�&��Xn*e̐ӏD[Ѵ]�-�fu!��F���
O��~o/�OA'��IT��ͨ�&����[�©?dn�cǼ�=-����}�"���a�=�������	�hs��WT׭K�n�m�-,���p���H�b1���I��T�>Q�D��4'��̴�����ISq+7[��4��<{�Z�-��:��v�(��2^l�rm��5�^� yl�$�����'��Qz��-V7V)�6�8���� v"�m�)"�3j��/o�S��'n-)�	V��C�Hǯ�e��I\��ƚ�ȇ�2�2q�|��r�3R0��a��C���=��8���6\b�SSV���}�Ph(CС�O\D뜛̄��̏K�c��kŴ�Vm�]�ծ���?��twb��eF��ҽ;��&��Do��L�{�����m2��O���ƫ/AΓ�7�=Ԭ����*��Τ��x�S4Cw�[�Z������S!�ף�d*Y�-���/�9%U�y�f/�ʗ$A�yl��a��Ֆ:���%�As��v���͋嚑�g	hI�0܍p�2+�Lk��	�}��Q�_��lh5@�P�3��[7pw����)"H/�z읲��xQU:����{�k[�\}M���%�R_b[yA�g���C��G�Z���G-�Z�g#�A��F	���L$�FP�A�8�mk��3������>8�^L2�~̭LŨ��ʾs��wUk�ww���9��dZ��!�}Wh��˽-�;�8%�a�VrPJ�@��^��a�Bd��W3�8F�b,��b��~��)@m3����~tkk�%F�䥗}��
�	~��Š��RmYс�2�8D�Y���
��!t������ ±�%{s�`�I���A��(Q[!^��"A���u���������MI)Ƣ�,a��F{`� ٪���|��2�ÛI7"�s� �Xl�>7��MV�sx��%��U��Ȱ4֥><��#���X%E�l�I*@���/��:���O|���S�p9��^�<5� � ��>]C0[����O)Y�9�S��P���V�x�OAA+T��A���H�i]�� ��۬���.�/��s!"O?�K5pF���N�������};����ֽ7���@t��Yt:qۣ~oy��sο0=��Jⶽ�݈Dc��g��f�H�~������a�'軆Ԥ�������z`䷈*gA墾]�^��!��wP���áb/��E#�>������h3֓�ρ'���J��UMF�	(	ҥ��������m�t�8�e���"�%tӠꊌ獙QaVxç��[A���|( O,�l������S:ظ�2S�aAw�_�q['Yx	�6��{�p2, K����0��5�`�}�y�D�?J�09�t X��8u��&�+�m�Υ}T�@���_���1�mZ�|�mǀ2P�T�3�w/C�e���x���'�s:E�P:g��bC0��n��9>R�l�$R!bBW�*��+Jr���Y��x�'�/%c{���R����.|1
Sp�̎�h	�Λ(��ڿ��<Jx��p��4�a7�(C^R��~�*���@��݌��ax/��}�d������=Vz��e�'�\���;��>hd0��"��2���u=b�âsۤ��2,矬�/����0��V$$tu�#�&V'�5�E��w���xGR�]�����_������f9���,V�g���4Gf�0�Ŵ�FfP�Ȧ����Yy��~���Ua�y�bH�������L5{U�"�1:��E�\O펆@FK��ȥ���U��,�^�ʃ�챻!Te�h��^蝞o�U�	�B�ѓ���r{��"�|U2�Vp��(ܠ�ON7�[r��N|�E?\?�O�,��g5؅.�����w�b� �j$J��g�a�)�ר�<Q?>Ry���B������rʱsB:�c.����(x�N�d�H���Ǎ�?5�U�_h-���E�B��1i�9b���S�< �:踪�����������ڍxG⑀��ٜ�0;��U *|C��6)�B�D�o̦���.�W�r��$������������5�Nd.�e�,�A�V���nr�s�<����5�gxf��T���'Ռ
�?E��p����*��3g.��(,t�0�D�Aa��ILl�����-��^!��BXy5*-�m��6z�ˆ���>��8Ǚ�3��t{��<�Z��.=D�+��?� �JIȤ�"㷥�E�D��G�n����Ev؏�Ŕ���ڃ�I_��zN����?�|��F:JH��Sf<�5mT[�+�	b)��ʰ�8��'��z9Ա"d�N|ͭ��U���N�V�j�O'�Yc�@|5w�Ϡ�{��,dkl�Owζ�U-�����38P�i��mp�?
�5�^��8�G�BFJ�Qoz�;�j���3�OBښ��&5D�A�,5����Z���Vh��������xmo��	-�L�����]��G��m%�/DeL�k��^mO���π0
��)��O�cե��~E�,s�G��f�C�D�Ner��.�QZ�$m��,ʹ�X �e�ἅ�p���N�v���f���G���8�T10�ՠ�������k����0ΐA����ø�j�i5	�O�9�/ e��Q��!���������缩�Q��qj�ܚ-v���j8[�[;�cĬ\v�Iݪ�WKt�԰~���Lsj�H�4��{���'����M��W�޷��>��M�E�'S�!B<S�%����BCS�������Ӳ�~��ŏ���++�l��S�����.��X ]j�����q�ĶJ�gV��38������T+�N�\�+M�_�>�`7?JG�����[M�����ڷ,��2�4�k��?@#l����G[�ֵ�o�ҭʭ5���;`��@��V�o�֒@�X6˿/r�:��o���~0k�TU�&�2�;�)�k��$lzY�Ϯ��F��Ű��G�Me(��y����Q�܏��7�te�''L�;�-�HW
|�&�>WX���~�9����k���L��_��b��O+2�A
y3L��$еp'��ٌh���Fx���P*ߓb���R��h���4x_�����7t�͂r��
�������%)�Z<�3�@�.h��hD�i��泌�c#�����nvϥN��/�i+%����GE�tͿx��tc�{zg+TML��s��,ǤLᵨ��r�M�yШ�7M�[&����*��1�W�5.a�H��W˾:'�'��=�B��w��t�����H���x��wn85��s0<�~� iD nm�q��O]Eu�$�%�mOX5,,������6�%�Jv���T�G�/�/>�o��<5{Tz���GY:X��A
��V�f��9 cQ�LH�ԩ���Pk]�AKv[���]��lp>�J��[�6��R;����j	�ҩZ^m�Ϸ�Y�q3��Lg�ۺ������F��Pjp�:G��<�ȡB�Z�Io��e�_5��q����vC���+'��$�t7H���J̱qDL5�#č6b�"�h���e�q'� OL閷!t��>�hg}`�1O�+�	ҏ��5kJ0M�Yod���gs�+�rvgb�tk��J���Zl��{�f��?������]I�����Y�����d�-Z� �=Q*̾K�Q2�wW�7ծ#܈��� Te{A���0���ͼ||����D]�j1�	c�E�vd���Jfۢ+_��}{��%
U}��_bc#�8<)7Ŗ2��P����!l3�>���.c��mjA�w �m��l�Hx0������bnV�X(�9~T�d�(��N��
Ϛ��}��;a�F��%����q!_��8A�7�p�c'�_B���aw��@�8�	5*�O>��we���c��;�#�2f�,�2\> �����m�]C��$p{�k<62xeT�0�u3�=�x��R붣��U�m��ծ:�o��3�1P�,����	[<��D���*�� ��P~X����A��?�����U��u��f��8_�D��P��b��k_��t22	ذ�N��P�����9��*�I�Pb���]R��B��8���_:�$�Ǖ+�E���aMZ	�Z��� ̫����9�d��7�q�zq�̹l�1p������0#��������3c�z�k=��*RL9}3H�?��IԽ4�#��]����!�*n&���m}�[��7:�:��N}G�=�JQ&�"J��������\����j�@���f��rp�j���P$����5���bF+�[�s��z~R�0�g��]2���U^`3�4�o��(��_h��훳)C�!���0L��g��;`�x�3��{�����a �;��m(x���@���1(�O�#�]@����QuZ�0ב���'��g @ϐ]{�l��N��������fW4�p�6N F�z�]O}����E-�-;C)��q^@A��N����*q���t�zY��7~�E��3�`{�#M��Y��l�Ǹ��,��Y�6I�����lb��:A����O��>g�&����L��^:�c�M���n�F��{�Ėd���״�]���.;�� �Yμ�'2]�}C|L����"M�N�_��`�l[���X��$ix
�m�t���\�����M�3��,9+���q�]��*��8{��/�*J�W��.K��r{?�ϳϳ�J���Y�zI������î�v�GGYzfU=o��)d�&P�� ��"#{PT�*[�5.����j����c[^�2(���*|�diǀ�J8��3��2�ӧ�	��E�.6����CRf;�[{ 7�?��$���'Z\v�]`���TB�~�W�l��+��2���s6��,�<5�� �?�[��̜�,��L��(S^�j��&%��k߼�%�x� �����۷��^�7��L/��
{�t��o%a`����lN`Gܫ#%��1��o[9+�Yj�X�K�N�C�c7������&�m�~vi�m펕�W�p�81�>��I�@2j�$��J�n�`S�;x����$��Ⲡ�Ƃm+��a��X$�ı�ä]`�BlL��M"���Ёv��4����RK56���%kQ��#����~�b���巘>�Ǉ�HCM	E�«�I�)<��
���\�W���֑	�c�+1G�CI�,���/�JFTȵX�B����Ƅ�Z�_J�V_�a8E�f��3�0���-,|��Pf���غ�G8s��|���ط��ڡ!��`����=Ҝ��e#'�,[�A� �6�0�,Uq1��}=�ZPh�/,s�9�2a��wfW�ϝ����z�Z�7_�]�T��b�6ɑ¢�R��a�Z�!c �yt���p�o�mN�����>N��,$g��ݓ2�8fM�3}�6��[�0���`�[�Χ��LG�o7W*9Gb>��mp#6-��jobS7��̎B�N��	�aFQ�3�d^MM׭Uu�j�*����\��D|�����"Nx2�FrX9<�j�!��B{������Y��>�?�u���a��Z��"C4h��A��P1���/��c	������s���X�6�ӂ�ܳ����fvPg)=����d��u�4�ᦀߊ>P� SPS��P�nM]�H1��gia�C�ryA=����7�jUS�;�Н/��aZ���#s��eȘ|K��9ME���^b_��OAV��6bǟy6�U���X��5t+4!�'�v�3�2P�*�J���|sia�ơ�l��z���"sE[3Z[F3 W��;2�t���pj�8�!�Ui9���`<���u��5��̋#�uld��k�b��ˁ��u?�2@��ޥ{q�����jX�c��T<g	�G���&@��0��GW��W98F���gk��F���M�o����M���8�J��1Dp��+nhB+s�8y�8G���_���t�V,0�?cQ=)����e�Y�v�%���S��>�K�_���,gi��XK�8S������%������&B�f�%Q���*%��ꫢ/��q�("�s��O|S)_���j7/�]a�=tQ]I�L�B2#��%�s�� ����]c���G��Y�

�Oy�F�5��S���ֵش��o�N,3|�O�:��?�b����e%ˬ��s��s`���{g�T:��Җ¹�Z��3�_{,jk��_�Tv�Ҕ�k�zD�2�wx5��>���
6J%��#h,/�O�I��]v�i���9�U��'�Ꝃ��N�?��NF���Y����"�>�$�%�u��Z�k�LRh涄IsltB�J��T�[j�JY��aG������GĠ�J/��#!� =�堂�ф����Y����LK�ve�!3�;	�QVX}�9��5��[F�|=���g��+��� �9?^S��B���T67R&lE�֣֖�Gv즼�,�]�.9�����s��M�"�nGY㮻5��Fo��c��N�	�O(M�x1�Ϫ���y���3&���J�K���^H��A�ಒ] 0��i�F!�f1�������Ń�+�sV-e�v����]v/�g ��B|+�yk�.�X�M����7���7!"h���W�;�)U�B��9�n�^��u��Y�gX�����]e����:����5zuRuy�'�Y	��QK[�0������S����K)�(f�����8YlGJ8�[m�Y�r>�/��
d��n'�NLk�n�:���ę���J}n���2!1'#���M=^�S[��3q��Qɱ7ND����Jj�~v��N���%�.�:�����>j��מ���iY��_�,JZ{���=/:by़�R�`�<�	YڲU+g�5�S��a#J:���v��u����8bc�h���b6��~���Ģ�7j���r�U����TK�1_�[�{�0��B�z쮊8lJ*y�?��6F=���ָ�.�ق��^ ��g����\gL�֒XԔ}f��g�`sc���z3驍.f��uS��I�����ȣ�����40�,����p�e�4����o�8��M��pO����b��H?���=��N���CI�i�lm|��	�A����Y$ ��9ֹ�O��&��C��.�$u�i����W1��1ӎ���'�������+/��-��g%2d������Y��B|ꠦ3!���%�ظ-~3�rأ6ǯ��$��a�*�><�Z���Pwa1��~`�����V?X���dI�@�r�^�NSotaO�����#�nD�$v:���w�d_���L��3�Е�C)	;;��0��0�=�GEI�8�0`j+�y�M8�U%��R'U�D^1g̓�X8/�P���H�w����7��a�Ry}Gz՛7�z�`d��qq�j���y��d�ZO����a�.��r�K������f�)��N����	T_d��V1��v��o�XEU0�a�غw�k����/uI�+���x5XM�s���5�ǁ�t/D�.߽��S9 �iP�f�}H*-�'ʮa�Nz
,;8޴F01��!Г�H���MV���<�Ox�	�z�� 4<\o��澒_��b�x9�&hg+�4���?��+����	5]�j5]�&��Qwi��*Ql���~����ίe��<Z��Ӥy�2VV}��y���o�(Bqp��9��`�x�
��f�����	�m��t#J����Nm��fJ5�Yk׃ж6�����7���;���5��^C�y+��*V���1!�Wk'�p:�sM2�7�il��u�=#&�ϗ~Ut��>�wxϡ�{�=�?.���u���ob���[����,���a��L5JZ���us�U���:�{�&^أ��l�o�s�$���Q	�����E�}����'V�o�X@���?�͉��I2���&�U�{���n*ǟ������ ���#&w� ?��Xߧ�� �J-0Ȝ��貵������p���ԉEM��TzP��e6ӭ���g��c����޵�m'QBq��!B�:���c�чڢ�P��{�!��'���LcÂ�c�����IJ���o%YdQ��u�~^��VN�0d�P	�������D�8�O����k�n�����~,'����������
�謩���0D����3����d��B���d�0�U/�p���0iYB
00AL��4x��:D��$]��!��O��Q�5���@��f�����5�?��"�<+����.ߘ�>gV>j��Ԇ�r��2>C,ݤĽ��S��/>�k�Q���5]�4^�
Rj��n�v@2P�����hd�My�b�Q��Yؕ0������Ӫ�+���vߋ��K)J3�!�eޗ�Ɉ��Le����mpT�b��/炉ӡ�ԭ8}�v�j$Wo�]kΈ|���W��ys�GФ��+h��ݯd��hw5#��$���EB!��=XB<�Cr�/�iD(ߒ�?w�Ө��K�L�W�;Y�+��Z��~���4{ܩ�x>��x����t#�������B�^��4�9�;+GS�ǌ���>��RX�@�\�L�������HӢ�������L���.e�a!F6!M|dG��[�N�\��Aq���׊�O���ϸ�=Sy5�z��kId�i��X@*-+k�P ��XS�RB^a�8����L�L� +w����1�nx��e���N�G�o�]	F�����+���<������Ϋ�4o|s"ΑÄ�d�F>���8ĞVc�lC�PՋ1z�E���=d7���!���+ݲ�Yns��l�9��gꈩ����]Q�j��N�=ex*��]�ƶ����憪�p�2<=�݌�P6{�v���� &���D���F���?����ܬ�A�A����_�f�03a��O'���Ә�� &�r��n�we�vC�
�H�bӹ�O���E��HSgbЊ�M�Du������,2�J��&&�#G(�gz� 
`� FB��)8��7�)3~.<�hʘ�z��j�0��Ik��ƌY��F�#�x8~������-�Ӈl�,���G+�́�2��>ɒ�9���:F����9n���K�������yf��>,`��hr�[ 쁕d�26��,��}�#*6=���L �ر��^�?}8���2sRf�~^a]B���'8{X�[�uI3sT�/��u�!䁯$%9�w�v��pOO�{Ő�hq�<��#,%�-�c�_*���"���I����Zӵqdm��c��z�z#
 ���p��y�&E�#F�r�&��k����/����-��s�ف�.�:׹�zl�ݒ�%�ń��x;,�h�7���3A�s�/l!^<�`��C�����
㞹*{�%e�`�wur���f��,5�+�@���Q�w�b+=? v�o�3��	*W���|bMAO�G|g�G2���$�%f{E���e����@Q���`����<�q��)�3.%P�Ӻ�K�� :�zz�հ�EjB�8�7����_q�P��l��=���Tn���N�R���!�^�1�9�����4G ��9���.�UV4%�@���噜&jV��#�Jt,������-��!��~���m�F,[e�(�I��u�;Ȉ!��P�~�d(OGk�J�ʹ~�G(Y��a�,.]����B�T�Y�v�o�w�>�C0"��JL ���zv��d��g�
H��Ag�I=��l�"�Vd^fջ�b��e��J�h+��;�]�@c�m�S╘Vz;`T"�!u�ώ�.�:��Mϸo	�t)�POe��ʅD���n�Ҿ%�*�����W�O�C�V3��ţ���TЗ�N
y��Ć�G������WlZ�?��m�ҹ'�O��-x�������:.)��9�]M�;�0(yȬw��9��@M�u�ݺ7��U�����R�W�U�����~.�W��C�V�'�
�H}�N����^�nƨr��g[j��l�\��hN&��i`'y���g�J�cF�p����d�����6��8K�A�y��J?�0�圥o��������j~B���g�;�����ߵ�S$5��6�Uw�A9t��H�A9k�UL�`TV�j,��a�q���1T�V��+�ܫ���^�2�9B9�Z�5ݝ��U��!���6����(x�$0�
���-���`\/����!��I�!Ϙ��\�q @�W���ޣ��d>�u��)G�!��G��O�ׂI��]�UZ��3�����?�Z���(v��NN� ni]r?�g��[����]rQ���f��Є�'p;����Aa����	�5Z��	߀M	~�&S��>�V�V*�q�CaJ<���^�gB;��ғ1@Ί_�P�v�}+zp�ʐ���(��J�b�\2	�1j��1��=�?r�0���w��IJv��-,�ėM���?�����-D�̮9�>�o2/\U��ք.���"LLL�����*'���w�����Eؿ�w)C��{��M ��E�H��W�4Ot}����1�*�^wvӏ���c�g���7�8G�z�ːj�D-�*�`u�� @��C���H��Ԏ��Ԗ�������6���<y�1�ɨ�r���%a���u��<��%���gODV�3�}��x	�l�o+��P�r�}c��>� �=���R�&����Ӽ�\D)��l(�b��U �����B��`���u�BV�ʓ�:�\�q^��;�r���W��q��@D�����Ub�G�� *��Ϥ�.t��d�+)�����ed�����PMr��fp	���c0��uk49�\<,-�:����u��Α}�p�Z�B��k��xO�� x�mO$���&%Shv?�����T�Pf���
�C�]��jb���q�7��o�F ,�B�/�uƒ��$(�V�)��!�I��VR4=K��=,M]+g�g?Π@�1�Pbv\>�$v����*ί�KV��6w�r��x���R.��QM�6%⎍n@�T*��.�w��r�.Q�0읚Θ��}5;!,ڶn܂/[@�r����DXƃ����&�?4�	�Yϯ�4A��U9)�]=abV��"�
K/�5��"��OX�L.8�o����׸-7�����?���1�AE)�з��^���E���3�	���d�Ɏ�oгk�'7���|q
�'� ��D��k���
(�̗�����8g!��U-�tV�pqXg�X�m<��3޾�n�9�쁉Y
��������)]��R�_����.�˅���`�a"�[\��Y�����%^���6�܏桂��������ͥ�,�V�R�AĂku�E���`  �K��ڛ�N��[��9��+Z<�0���P�aA)J���_E~�0�AR���Ä�@�	V���ŗ���QQ��������/�*���E�n�8KZ(��z����je�4��[hQ$Z��/��x�k;���w4fñ. %a;J��@K�Z9�ӣ���s^⾨|�ׇ����?��O??��B�~�0b����K��3��qO�����KЪ.�u7i(j��x��]U`�:]�\��t���7v�����St��KےaO��<>�`z_Ca֯�T��h/�8�7ZS����,w���u���C��H^ǈ>#hf��a^欞���᭺��o=S���� Տ0���y�0|]���2��O@¢��@N���� �Eյ�U��I�g�DG��*��o�-J�x28�F�?��������4�kg$M$J�}]�r�p4dN1*C�yPb�^^4$���V:aO�o���>H������2��fr����Λ�_�]w�����ןvev`��T]�"C��y)	x�����e���'��PɝY���9A��Q!�/�h�B�8���i�c�����Ũ��R�#�nD�[ǆ�0wCIdcjЯ�f�j	e�O��j���-Cl����H�MR>�1��7d��:�D�i����PH7l�l��d��W��"G�l�L�M­*���s^�`��u��i}�ŧD��ۦ䅜�t>���8ax1os@��n�؉@zqwjX��d%X��N=��������F�|����N�*h�~mt��^���J9���s����!ȉ�#�0�����mZ�AH����!��_{ |�,�-ߜ����N+l'�'<Cz���(�*%�d�VM[l���Q���_�C�S���~�.S��
�!�=�;��[�9�;l�"�5��7w���Ղ���s|X;Ņ�����Ş�A��SwaW�������ѝ�L�N�#��̃� �F!��PU[��#~�[+>�P`�{��z�dײ�rX�E�W�E�<�*oH�xL-_K���=J�	C��׆��3��cP~�@�%��v����m�9�4nSj�����0K����Y:{`X��{��@o��[���T3�A��fo���$B�m4|�w?�_
��iH�$���M�4Ӷ W�S��3m,K�c�$k����Z�p����H�&�#(��ڽ��Rh#���Q���Y���ǿV1����$�k����}��=�6�����.̧���	��\0s�:�;����,��!� !*!�!��Vg��~�����qV���PVTMme����d���m��D[�;��u��O��'!�$�O�	i8G~��y�����~�`������H���ޞ����I���U���HZ�Y�<ȸ�8����?��=�i��;�n��'b�m�Du��v50s|!���?��4,��B1�Kժ[j8곫ɴ�#3��zT�/V��0t*�'X���9�R1O��h5ab�6ߞDX[��n�����ۤg�y+�_֌�r�K�hMA�����]Q�������7c�;/w��}<�Q���?<_�������V�'5=�-�A����T}çS���S�ZC�?�B5��ߪ�?�|��<�\��K�l��^j�dt 붕# �i'X�ҩ��T�Xd���>p��x�6h�L,7=I[�w�RzW>|��lTV�t��D��|�8 ��� ���3���;�r�LO#�\�uZ>��5Dg`;�=�k�э}�i@�����N�Nc���#g#���QK]�i<�vS9T��.<����J��d���X��w�8avh��aoZ�aT�V��Ai_�Q����M�k�̃M����0�U�5��Љwߧ��Z�a�� d�e����u�6x���*��ੁt6�{�I�p�xW���,d��d�e��l&���>�''���d���z�N̡�{����#���J�l۾ ؛$�b2�Q%U����h�/�"�=�
�lG.��f~��J����}�)qbMF���6p�=WUŉ�t�
DX�D�ƙ�pZ��|m���V%��q�鍂��醘= ��H:�)�@�,�O ���R���?q`n��)�|ӝ�p���I�f�x�k�n+�MȒSPQ�*�ʅȌ�ҏ����RU�YF�BM�˄�$ߩ�����'5���j��:��Ly���oeu�3�Ky� tE*��� ���U�d�J�c�;�L�T�C�a�Ȝ������ � ��Q���Wy�h[v2�/��� Z'^���R"�l#3��l�ІY�H�2���<I�@~��,p���K���_'�3w��v����+1��6;b����il��F�\,��������9��N/��|�m����-��.�꠭=T��b�~�u�G=顭Q�C�%�»0Z����1�� y�'(oj"���[��"Bf�U��^���9����zC�:�&HA��T#���?�6�ݡa�!&)�k?��v �t?r���,$���i�khd$;h=��Vޔl2��z�?���.��0��k,�+�ϕ���g9m���uX��������*����Z�׬��[5&�!�GIsi|��hnGJ����=�T��U��T���c��}y�^w�Q���@J_{&�b/��b�!V2I�@\`�l?��vJ����/K�H��Ud�P��As��ۥy��r�i�\��6y2��ڍ֓5����
�_�"�ڂX��O�o`�������;�,�1
�U�'ԉp�x`@�"y/���4�=*^1ϔ�F#��a�j�)ZK�����<�9��IYf /������Q�૓D	�&����D�.?mc���TD�*X0߶)����� �����D�$��/�����?dTwu�[Dӥ`QA���[5p��.y��҂�;�iG��Ea&E�o�.ǹ<�� �[�0_��M�{�]�����YBOK@��wǽ@`�w5ZtԄ<��
i�5�=��)/��%'u�0ͅ&i�;a'!F��V��Siͧ�.�w؎�ϫ���5���������b G����jͲ����ᚓ^'A�Vr��B��>���z�P��%ڷ��J|k$<��ִ�_�<���b/~����`G����B��M8��cW��f��Gk��,S�@��>'[>9y�v�^����١���N������#�� �H�򀇴*b^�x��(�w��Z��	=g;���&%U�B[�u�Ѐ��Ƈ�p�ŔSo�
A q��ǵ!�LM���X=5"3�$��L�߃� �|F5�w��� �Qy��cG*����.�02��w$JZ¯g%�6�~D�s��7�콕���0˒dc�hx�ghs���^���x�_�T����F�ݓ"VRW?`�����g��u�~8�`��y��4��V�P�t�hy3nD^��>�P��M���f��V}(�^R������x��C�<�"v�Ӄ��!*��0U�
���ƶ|t�<�I����*L1���k�xS䩵"<�kk���(i!Hw5��-��2���k �h��9��,w<���<�1�Y�Ev��Hf��_�G��H��,�{�V{7.W e��U/�J�<Z����º�r/,Z��pn��X1���15`#�3��ֆ-زڢ��_=_�P��^�@�>v�u�q��o��*@`0j���kw����%��FY��r�����BC'&`53p���M%�_A��>�����������줘@���
�j�����L��z�Q2 ��ܪ��+�J��
:3F�aOՎ)���5�?�h�c�P��<�8�W�T�VQ�f:�azC������yx�Ԃ|���^$���Vn11^nI�'����4��u���͂L�ȇ"V�R}/8�$�������O_�eM��˰{��e�.N'������tp�8�&�6�� ��٪b��������E9�j`_���J[Mn�Աv,��k��^���y�Nü��y0�Id�u�u�\,}�j��X:�f�o.�٤Y���Q��Q&PW�֦�d(̧8+5}���j���
���w�UH�аW�P��]qoHvw���g(��	���5�~��>;� E�r��}���Y�m�E�R�>�?�-�d�ٴ�g4g�_CC�2�Y�J��(��S�́6--Y�uN$�+g�`p2@~�>�(���c*V��#��]1D:��yD��uu��Вj����9N\�cͷ�@�$�*g� �xɹ��S=�^3��|���Fg��֖�g�7CÉ���R���y
:	E���"�YLV}�qY	}�*
�v�56���HF��Y�AG�ɯi�l�E6ښ�3:�Ro8�M�RmN�^2	 9��pG`{Ԋ���;-������M�q8]���D�s핵��8��D���s�c*��[������ףW�h�T`Ⲥ�8�{�f)'n����{}�-�ެׂq\�&&I����'��Pp�b�9	
S�^K.6�A���{VZ����4�^�"�O�i���x�N�2걷K0 4~�fߟy��a�".��wPu�l1u�8	h�ܤi��PrUE6��v|,?�q��7=�c��X�� ��zLp7�����>�A4TJfAU��g{qjp1;�,.�0#�fcӀ�\������w��Զy�U<�x��s[���UvH�����湌���b�B�t,6��3e�L|�b�X)R2�% �R�i�$#�"����w#c��C����bf�|q���m�]��Eg"\(�x��F�Ʉ.�� ����ھ+q���T��q��8�|B '��`;,e����v��8t�Q�i�[f�V�λ��I�ٕ:լ~朸LK�Nmǐ<ڟX���Yn2e�j7��,Ӷi����d�,V���HIs�QA��F���7%�#�����x���b�a��7��$-.�r.��M;v��Zy�Y��b	��H`� V)[�B<�T	
=��2�����z:�:��L'en3��..���-m]dv�p��^�0�=��`sa��(+��s?@�:e>���Z��ܩ���%��)�lk��`�^tK^�KGt<4�W ��$�ٮ=Vx�+^�mo�9�y5k��y|R�Yy+G�x,�q-�64I��+��-���p�_ �@�a�x�8��p�<���p �M��.��L�^��QG�~ $lI��j�o�X�A����ț�i4��l�ή�n\Ut2*����i<f��ı�{�o� �euOD��A�]Jt#|0����ty2��}ĸ���9�r�&A�
��b�Fj������8i�뻧��}�F
C�Y�����i���`d�T�Cf�.�i-��Zì���������~���TD?��4O`�{I\��{v.�gp�i�l��s�*�D�vȧtz�7�(����m ���>l�ֹ3y��p���Gv�a�j7y�#��n��'�py�-(%��a7�D�e�|_�2��=[�{Ӂu��
e
�pOT/(4M��S���J�
�=�/[s��>U�MY�k�M�6�9ʀݚ����NØ�1U�(�P��t�\}��F8�k,�:=��Z���	�`BY��t�T �(N�ҕ_�yǐN��At�G����q�>�&�mjvV�M}	����ɦV ����BhaV��C�<�W5�!��H�m��ܳ����4qt��8��s�Ls��䙆z�Qw���*_E�����	|�i�����D�~L>���:jT����V�E3LMa�͎,�,18�$���q�$ I��-8o1ae���x�d3������Rbe����6� ��]���/����-!����UPS�h'���H�������@5
�e�p�;��깼�7�zk���h;SG)L�ܦ�.Zjrx0�r���=�����gC)��2���1��9ҡl��._��������I��YF0�<�ސ�j�~o�r	jD&���`[!�#��D���5|�I� �����'�D��/��p���r4�5�d�خ��<�t�mv�)������h�`2��g�-}�ȯ 	�U�ќ��3}�<���{`�B?v�T�]_̀����nջ��m"���r��X�g�r�`�Q�[��@��                   0  �
   P  �   x  �e   �  �                  �  �   �  �               h   �  �i   �  �j    �               e   ( �               f   @ �g   X �                   p                     �                     �                     �                     �                     �                     �                     �   h          �� �          �a k          `u           pz �          (� "           P� �          � �          � � �      SeFFF~~~->�^��5�k �� ������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ,    � �  � H����*\Ȱ�Ç#J�H��ŋ3^�q���B���Q�ɓ(S����@�0c��)��ʛ8s��#�?,`���ϣ4G"8`�ӧPSpy&Q�X�j�4�ׯ`�	�гW�n��kطpwR�	ThڬZ�.�ڶiܿ�3H��ݪj�Rm��@�ǐ!�5[�(̟u�*uٸq�ϠN�|�pٲk�v���`�uѾ������6[��zf᪦5o��z����+���Ÿ�,y�z�ѳ/֞x���	
�H @���R�"�;Tx���	 _^�_��-by56f����|��g_N�w_~����e����^2V���G�J	&�@}ƕV15wVwޱ݅f��u���g^�a��\e�%!t��'�|j���G(��3�H��8�5�i$ZE"�)r6 ����O�G�@q�a�h:I�Q><"�܄A�h��_��a�{��'�a���N:�E�P���+��b���!�}�i)�5�7�W�YyU���V��\މ'�N^�*�z��iT؅��w�.����e��I�檫N
�Nz{'ֺ訞����
l���T���*������G�������֪��K�r��w������[������\o��e�Z���")�3Vzo��޸/N���v�-dnC>j�x�"�0��>��~�����2[�'���:��+M�ެro��g$����
�K3Ky������<�@��I/�B�����!au׎4/ ,�<��{�\.�3k}��%[U�es
Lj�E~��V����os��(g�,�P?�$��}�����܇��.����(�S��Г&y��/��Q����R�Z��W�<zF�U�o~!�f/�:�V'����'q{����B
���{?��XM<D�����t�<vٽ��x�1�{=F�Z���ݎ@�^jX�������W+c�ْG y�������~k��,�-1eL	iI[׼���H�B����Jd4���B���,|���>W>�y0"@������wg[!��ת�! tKJ�jX����e��a���C��� (@@EHQ�"$�RN��<EO�lU����hL��XE)�h$<!�E��.Sd�Hϸ�>6��U��A ����[�̗�%M��kd���6Zъ`
��8;��TH Y�?�Q�}$%��A����C[��P2����#*S�JVNэoD�t0�X��a(GyI*��إ���6�R����AԻb�(v�t�-��@:3����9�M7
��K����q&���D����K`�3�b�U�w�K���$'.�FiNӔ��5�9B�QU��O!*���ѡϤd/��Nwj�>A���
T&�*����>#j��Lc$7�W>mԥ)'C��j
ҍ%զ�6An�ɠ�k)P��\������:'
L%� G����S��o��P�R�5�IUj��j0e�h<vm$LUyʬ��\�k��V$)�IPL�V ,��l-�V[כj�K�a �f<1�	c�:J\�R��d%&��կ��H b�֡���D���c���Ҕ�6����*��j(	��lY&����h^c�z�ަS���gA���/�����x�;ک����e�[})Q�:�Htլ|��\������mnK��Fӯ�|dpK6��O�Mn}�����7���o[!:YlfW��5�����߷�@�+z���~�@��|a�a7����iu��U�R���{]�$�h�.�oXc|^�bu��\ge1l؃ixð�	�����M7���o%�T;����2��keҊ��ZV�-;��X��	��s�fB�����/��׮��b������"�v��M/�Y)΁��c\՘���"l���^6�����;Kd�:ͪ]skU����Z���iO]bwY<M>�|A-�����E-��KE�.�Y�{r�]��Ђ���$eH/��
/Y�mv��~�fWٳ�5�����b�z �ݛY|[oߖ�},�S�h������qr7�ao��H5��Qc�w Hbu����Ŗ9��%&�֭^�N�u�>���P��$0���c���O��遲��p�����(g�b_Ü+����^?;�{,���hב�zǏ^w�{MpCX�RM>��*|߶]9˅(kNk���Z�ǣae���-ך��iR�P݂��u��s�`�NG��� �% p ��g����������7 �w��e� 7� �; 4m{��~\�r<����'B��/p��coy�8� ��n�tG���M�C������<����(�C½��@�~a��3��{������n��x k�夶��0y2�=����&�}���d�������^��'x��ڇw�y�Gy��s�Ez�w~/�7����x������'� ��x|�'��w�E|M{)�'8$���4��x��`��o�z�x�D'�)h���w��~MQ��7{�W�x�ф0�yׁƑ Wi�|�5�T�zIh��G���|1�)�}�t{�n'��d�����Y(.�6_ˆvc��T؄�g���wxqh�y��7y���(�W�=�y��!x[ܶ�iWhHq/h�~G�=��x�/�|O���h�v�#�̶t.vH�Gh��F��(R�y����(�g{E���H�GH,Ne�,U'��.�}hy��}�犘����7 ��Y.(C�W�yW}�8 ���7?�G�Wyη�}�?H��'��7����X��w�����o1�i*�T49:�8�y��{��y�8ɑ��	$	y��A���Y'9������� �/���$���<ٓ1��M�A�9IFDi�!�)BG	�B�O�D5�Q�3�?��5i���Ĕ3xI��K��X�7�S�C?9��@�j}�}R��y��Q�bٔb���іn�y	!�-ɗXْ&����w�咂	8��{~Y��)�X	����'���y=�'�|�ǘqwLI ~A��t}��{���)��i��	#=a��w��G�E��sY<��W���ؕ��X��	��9��I��Y��u�M�)Y{�7���w��+S��"����d���ٗ ��7���w�){�9�i�d��B��	�P���~ᧈ�y�,I�����Y��ɞ���"����`9��	y`٘ǉ�)����x�����X��)�$��/�yṟ+��U����2
�4���ٙ�9�_9����ĩ�b��.J�Bʒ8�����7�T���W�rȞ+󗘨�'�2Ċ JU��f�Y��kڥ0ʏ�Y�~��q���h��ɦm
�Cz�J���%)��)�z�^*�,�������������:�j:�zڣ�ʟ��Z��=�����ܗW**��ᡙʩDʡ��~ڧbʟY��*�����h�0��D��#:� ɨ{ʫ�:��|Z�r:�MA؉�0��(���J�	����ʧN砒	��z�@z�o���Z�.*�z�py���Ś�}���ڦb�w������̹���3h�	Ѯ���I����5���jy�z�oX�o9��*��l����Z{���s��
�����+��گ�)�oH�*�����b�����"���7�&+�1��ʱ�Z� z�ȹ��y�a��)��I���>+W�y@��B˧N��z����2��e��&
�
�
�?)(;��
�,����*+��J���6+��J�F����,��4��1ڡg������3�y���:��
�By��qwS�Z�����	�[���K�Aʵ�X��ۨ1��گ�*�W*��5��:�Uْ �������K�(K��ʠ�+������}�[��ɘ�;��۸t;����X�
���9��b���$��g;�����k�К�5�]�����k�h#��M�����ɾ
a�%;��ʫ����:�������)�A��к�}*�Vk��a��9���J���ϻ�̹�{�'�����񪼹�"|�yg��[�L�.�&ڶ)��Ɋ�X)B6��暿���h�����׉��˙1*�r�~�������l�/l�̼L�������̻�o�~<��ŚD�.���AH|� ��L��g	��Z����"kw#��!l��)ÊV:��;�䨾���������l�6���'������@������J�bQ�p(����L�Lq���YxF�y�z4�y}e�@��}��,�� ;     ~  � ggg���wwwGGGWWW���/?�_�                  !�NETSCAPE2.0   !� 
 ,    ~   � ��8�ͻ�`(0��l�p,�tm��0�e����pH,��% %�Шt:�Ԭv˕*خxL~�崚{��pd;N�������~�d_��]�&7�����5�:"����� � !� 
 ,   	  �ȉ�M8띭�S(F !� 
 ,   	  P�)������L`�I�8��p܅�,���LG !� 
 ,   	  "P�I�:8�=����d���Y�c�����{jE9�G !� 
 ,   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,$   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,,   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,4   	  4ȩ��؞�'�����'�����	�!ۚI�6Rɫ[q�T�C78[�9�L�1 !� 
 ,<   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,D   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,L   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,T   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,\   	  0ȩ��؞�'�����'�����	�!ۚ0(�n�q)YҨݦ��j���# !� 
 ,d   	  ȩ��XM�{ݒ灀ؑf�*G뎠�kjն !� 
 ,l   	  ȩ���^���݇�bTG���� ;     I  �     '''???GGGWWW___gggwww������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ,    I   �  0` �A� *Lx�Ç#J����D2F@�1�PIrb��4X	��Ƅ0(��M�'#�Dٲ��.U60� Q�P ��ʣM,��@�@��*Ř�`F<X �@P�>d�����n?��@ �ێ,�v�:Wcر �����r#x�K0�(��ِ�3Pa� �2#a��Mk@�J�|3`�8�
��ʚ�fӟ
И9$qΆY+�|w� w58�X�F�kђu8�8��]M��&@����V;���klj��^ ?�� #� �i�������AWݑEX]q� ~kq�_P���6�@�q��^+9�[�:	`i]9�҄:�hڃ $��[ ��g�!�ׄq�" ��e�l7Md�HKr' y)դM ;       (                @                      �    �  ��    � � �  �� ��� ��� ���       """ ))) UUU MMM BBB 999 �|� �PP � � ��� ��� ��� ��� 3   f   �   �    3  33  f3  �3  �3  �3   f  3f  ff  �f  �f  �f   �  3�  f�  ��  ̙  ��   �  3�  f�  ��  ��  ��  f�  ��  ��    3 3 3 f 3 � 3 � 3 � 3  33 333 f33 �33 �33 �33  f3 3f3 ff3 �f3 �f3 �f3  �3 3�3 f�3 ��3 ̙3 ��3  �3 3�3 f�3 ��3 ��3 ��3 3�3 f�3 ��3 ��3 ��3   f 3 f f f � f � f � f  3f 33f f3f �3f �3f �3f  ff 3ff fff �ff �ff  �f 3�f f�f ��f ̙f ��f  �f 3�f ��f ��f ��f  �f 3�f ��f ��f � � � �  �� �3� � � � �   � 33� f � �3� � �  f� 3f� f3� �f� �f� �3� 3�� f�� ��� ̙� ���  ̙ 3̙ f�f �̙ �̙ �̙  �� 3�� f̙ ��� ��� ���   � 3 � f � � � � �  3� 33� f3� �3� �3� �3�  f� 3f� ff� �f� �f� �f�  �� 3�� f�� ��� ̙� ���  �� 3�� f�� ��� ��� ���  �� 3�� f�� ��� ��� ��� 3 � f � � �  3� 33� f3� �3� �3� �3�  f� 3f� ff� �f� �f� �f�  �� 3�� f�� ��� ̙� ���  �� 3�� f�� ��� ��� ��� 3�� f�� ��� ��� �ff f�f ��f ff� �f� f�� � ! ___ www ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �    �  ��    � � �  �� ���                  �  �����      � ���     � � ���     � ��       �� �����     �� ������   ��      ���  �� �������� ������  �����ozR1ML��    ����o�zR1M��     ���o��zR1��       �oz��zR��       �oLLLLL��       ��������� �  �  �  �  �  �  �   �   �       �   �   �   �   �   �   (       @                              �    �  ��    � � �  �� ��� ��� ���       """ ))) UUU MMM BBB 999 �|� �PP � � ��� ��� ��� ��� 3   f   �   �    3  33  f3  �3  �3  �3   f  3f  ff  �f  �f  �f   �  3�  f�  ��  ̙  ��   �  3�  f�  ��  ��  ��  f�  ��  ��    3 3 3 f 3 � 3 � 3 � 3  33 333 f33 �33 �33 �33  f3 3f3 ff3 �f3 �f3 �f3  �3 3�3 f�3 ��3 ̙3 ��3  �3 3�3 f�3 ��3 ��3 ��3 3�3 f�3 ��3 ��3 ��3   f 3 f f f � f � f � f  3f 33f f3f �3f �3f �3f  ff 3ff fff �ff �ff  �f 3�f f�f ��f ̙f ��f  �f 3�f ��f ��f ��f  �f 3�f ��f ��f � � � �  �� �3� � � � �   � 33� f � �3� � �  f� 3f� f3� �f� �f� �3� 3�� f�� ��� ̙� ���  ̙ 3̙ f�f �̙ �̙ �̙  �� 3�� f̙ ��� ��� ���   � 3 � f � � � � �  3� 33� f3� �3� �3� �3�  f� 3f� ff� �f� �f� �f�  �� 3�� f�� ��� ̙� ���  �� 3�� f�� ��� ��� ���  �� 3�� f�� ��� ��� ��� 3 � f � � �  3� 33� f3� �3� �3� �3�  f� 3f� ff� �f� �f� �f�  �� 3�� f�� ��� ̙� ���  �� 3�� f�� ��� ��� ��� 3�� f�� ��� ��� �ff f�f ��f ff� �f� f�� � ! ___ www ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �    �  ��    � � �  �� ��� 














���CCC























�껻��X1CC










����




�����X10�C









�����
�

����X10���C








����
��
�����10����C








�����
���������0������C







����
�������

������C







�����
��꼼���



�����C







����
��꒒���



�����C







�����
�����XX

������C







�����
����XXRss������C







�����
����XXRsx�����C








�����
����XRRs�Ẻ���C



�����
�����RsxẺ����C



��


�����
����
��xẺ��CC������


�����
����
������������������


�����
����
������������������


�����
����

















�
�������
���
��

���������
��
����������������






�����
�
����







�����

���zz1111MMM��








�����
���^zz1111MM��









�����
�^�^zz1111M��














���^�^zz1111��














��^�^�^zz111��














��z^�^�^zz11��














��zz^�^�^zz1��














��zzz^�^��zz��














����














����������������















����������������

�������p ��  �  �  ?�  ?� `?� `?�  ?�  ?�  �  �   �   �   �   �   �     �  �  �  �  �� �� �� �� �� �� �� ��         h         �                   �     (       @         �                  	-*0S=i�w��v��d��}�������僨⃥����w��h��X}�W{�`��k��s��m��d��h��[|�Gl�Or�s��t�ބ�荼�%% 5"Bi�W�ψ��r��f��q��y�ۃ��r��Qq�9X�4K�6L|1Gw=R�C^�A_�Tu�Z~�Xz�Wz�_��r��h��u���卺핿�(-"&=cT��x��y��n��Y��Vx�0I�/y3K�2;g))G#*9-3P4:_0?p/N�b��j��i��`��m��w��j��w����掽��
!&#0?My�u��~��w��]��;X�7yHa�$'F&5V-N�m��u��i��a��o��~��m��o�ڀ�苷쓼�!(+'316]�q�䄮�z��My�1Y�3\�"C "")#'6]3O�n��l��a��b��p�ۀ��t��j�ր�擻�&')&--?d����|��h��T|�Iq�<�%$%%%-U2F�q��q��b��g��t����w��b���哵ꔾ�*!&	<o�ψ��y��[��Hq�Am�@b�4"$$!'B,Cum��`��`��n��v�܃�冫�f��z�㏵땾�$+	%JZ����z��m��V��Dn�W��]��'+H$##%23Iyi��[��m��q��x����整�j��u�㈶쒺�$*!( *=b��퉰�x��q��f��R|�Sy�Y��<S�$ *5Gpd��X�r��|�ކ�懪⑲�w��x����펹�%'(-+4V[{�o��t��y�냩�k��Ow�5_�\�0S�;Ht:)5De\��^��s��z�ᅪ䉫揮�~��|�㉳�,2_������Tx�{��v��o��v��y��l��T��Jt�Gk�Kl�C[�/Z
 $%!(1S_��d��y��|�㉭鑱쓵��|����펹�`t�t����n��}��i���∫ꂦ�|��x��u��p��f��b��L��2Kw"*0 "":\��n��u�׃�挮꒰钴ꅬ�{�݈�뇳�%az�n�Ѓ��|��q��y�ۊ�铴쇬恧�|��x��n��o��v��t��O��'+CM';*.b��o��r�߆�牮菱敵ꊰ�����ꎴ� ,5W���u��q�ډ�智엷�튨づ�|��y��r��s��m��dv�HI�0$*X:!C56h��k��x�㇬莳땷앳ꊮ�~�ߋ�폳�	6SzX�������씲퍯닮�{��r��v��j��k��p��Nr�1-L/&d81T9Ml��p��x�般菲ꙸ싮�v�׎��*Blj�Ȍ�㖴뎯���拪瀤�w��o��h��i��iz�^j�R^�Kq�JI�_2.\g�g��s�ـ�㏲ꚸ�얳쇬怬᏿�!;b}���勪熦ᅩ߄��{��p��g��^��e��Yk���ۉ��}��fY�=:gVq�K~�j��|�≯锹헺억蔱ꉨ冲����BR|���톩�}�ۃ�ې�႞�w��a��\|����7?tE@]p_zI.8Q?Pa��d��Sx�i��{�݄�疸휽喵ꅧㆲ����r������p��|�ߋ�����}��h��Wx�\~����NX�,!0THZj��O��c��Y~�n��}�搱阹떺ꗸ銫ゥ䊶���BSn����t��l��[i�Yh�r��~����q��FYE09>JETe��[��h��j��X}�o���撳뛹�딻腨玵���*,Gn�م�ㅡ�DY�<Cn/k����偮��lz�<93>b��V��f��j��a��_��t�������ꔼ튯郦哺����22IoZ�Ō��x��t��j��e����Қ�曵ژ��[S|3 Uq�Z��m��h��f��e��_��v�څ�뗹�鐳匫耣┿������(QDi�h�ѓ�ؒ��av�HRz_UbJ(2J31@,10'OUxb��g��n��f��_��f��_��x�߅�勲斸퓶ꁠ�{�ז����-=kn��u��q�Փ��[JMb8!e7,N3)L-0[* 5-7Z��U��i��g��f��c��_��g��v�߇�꒶�������t��{�֖�쑻ꐻ�}��x�������퍖�s]zlA0o@2dA7W94L3/L-*?'U_�W��m��y��u��f��c��b��m��z��s��x��v�փ�ٗ���������뀭����3?crt��n�vPNtF5xM8lG3e@2b?2V3)P/;.6]��Y��s��y��v��j��a��d��n��e��f�σ�ܖ��������������鎶�`74|RE~U<�XC~QDtJ=kE9dC3_>/Y8/L%IPi_��k��q��w��u��r��g��q�ʧ�爩י��������������������eY�]Q�ZH�UGRExO@qL>jF4^>3W72H%!Sg�b��u��t��y��r��m��e��i�Ǐ�Ԇ��t�ׄ�م�އ�ٛ����������|�ދcQ�^L�ZM�ZL�XG{SAvN<mG;cA4c<.O3,_x�e��j��w��y��o��i��]��c��g��v�܅���듲�������づ�`S�_Q�[M�\O�TI�TIxL?qG:hG7k@+U<:g��k��i��|��y��v��l��e��a��o�݆�ꈰ됶�ꔽꎰ옺���‡��aR�bQ�\O�ZN�WKREzNAsI=kH:lB/WAFf��o��q��|��{��s��j��e��f��m�׆�茱떾��놩鏯������x�݈��`S�aW�]O�[N�ZM�RA~QDwM@pO?sH3^JW_��x��w����{��k��e��b��f��h�Մ�璴�����ꏯ����s��b�ǒ��                                                                                                                                            �     (       @         �                  �����裏������������������������������������������������������������������������������������������������틋����������������������������������������������������������������������������������������               ������            ������������      ������   ���������������   ���������   ��񿿿      ���      ������      ������   ������      ���   ���������������   ���������      ������   ���      ���������      ���������      ���   ������   ������      ���������               ���}}}      ���������      ������         ������   ���         ���      ���������      ������      qqq      ���������      ���         ���������                     ���������      ������      ���   ������   ������      ������   ���         ������      ���������            ������               ��������㮮�         ������      ��������Ϣ��      ���������������������������������)))YYYzzz��������误������������������������������æ��������������������������������������{{{^^^������������aaa;;;�����������������������������������������������������������������ڏ�����������iii���rrr������cccAAA�����������������������Ŭ����������������������������ƣ��������������������������������������mmmQQQ�����������������դ��������������������������������������������������qqq@@@���������������qqqppp�����������󚚚���������������������������������������������������������qqq������KKK�����ʗ��zzzqqq�����������������������������������������������񱱱�����������������礤�WWWsss������jjj���������kkk���������������������������������������������������������������������kkk�����������ғ�����������|||�����������������������������������������������������������������쩩������������������ʤ�����xxx�����������������������������������������񮮮��������������������頠������������������������㠠������������������������������������������������������������������ꁁ������������������������寯������ͮ��������������������������������������������������������___��������������������������߈����Ω�������������������������������������������������𿿿SSS��������������������������������ظ����Ӟ�������������������������������������������������ا�����LLL���jjj��������������������������������ѷ�������������������������������������������򸸸������{{{���mmm��������������������������������¯�������������������������������������������é�������山���������������������������������������Ń�����������������������������������������uuu���������mmm��ˣ����������������������������������迿������������������������������������＼�������������yyy�����������������������������������������Ʊ�������������������������������������������������ٙ����������������������������������������������������������������������������������������������ȫ�����������������qqq��������������������˻�������������������������������������������������������ʯ��yyy�����������������������������颢���������������������������������𲲲��������������������Ĝ����������������������������������������������������������������������������������������������΍�������裣�������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                  �^����ˢ%�\@E�4�WDB��{X���J������WT�4΄����{����\����Hn5�W��0Xχ�Kt`B����Z�]��x�A�����i㌷���|�?�����ωL?����W&�JX����\�G��J�S<�W\����W������t,?���N@��W\�-��W������t�?�?��W���W�_J�<�W�߿W��BT<�W�s�?���W(eB!�e �P8�C@A��W��H�S<�Wҋ���H�<�W�TH=S���W�����U(�C�LE`+��D��>s$��D��C�V�^L��O'�"����"�������4`\D�@�W0ȁ`�^����℗���t�?��DD	�_���ڕ�G1����S<�WZ}�Z�����NLݒ6�W���WχD(?��Ճ�҉h\3�U�3�҃C����1o?W����ϋD,?�?��Wz�}���W�t(?��T�����i\��jC�]��>`#�8a1�Ax X���Wd3�An"�3c1�Br��X�BD��L���W�D�X�����W���D��v��H��G�WωlZRݪt	��A@�Ar1�C>J�߁�\M6�H�Ǌ/d�s��D�J��.��[|�?��WX�J�ۇ��&P@I��Wã�0���o`����W���W���W���W���W���W���W���W���W����0�}��W���������������*�{Zk�[
D���_J����+C(�+C+�+C0�+C�+C�I�Wτ�`�s��˪Oz(z�@��W���+e��)���?���WdD���Wϑ�(C�h���ߖ �O��ÒyL4Q+�@���WO��ߟ��`�0��2b{҉`�ҁؐ��X�@D���W���V���W�������W���W/�4`�t�f�Uš!U�>�����A@�Ar1�ނDX��J�ہ<h�r��'J�߃��A�p�4_ZDӀ���[,B���3�/�TX�������W�OWEL����W"�Y�� WE��D�W���"�T�����O@&��W/�TX�����k�W�OWEL����W"�VY�� ݡD�����T��W�`����_J�׉hZL��LBG؁�`L��P�(�W�_����_J�׉hZL��LBG؁�`L��P��W�_���ᕈ��� �W�_B؁�_�� 0���_������R��ڸ�I1���\ �yX�5]ّ�8XϽ�W���'Ỳ=�����/�Y�������µӇ���@[mǈ� ����] ��@�L˦D���\�VJwZN�����P�x���H(������WX܀=�'��=�4��H5��Ĉ�(��H%��À��툜(����] ��B�\À�N4 /�����X��L�������WRǾ@s�WzH4L1ȁ\�SH=00�LiV�t�����W$���Z|��D� ��[� �eY��Gtކ�^��4B1ȁ`�SH=0�4d�t�?���W[t��LJ��/�����Z�It݈�]W���Rߴ����vI491ȁh�^�X����P좓�#��.�WωdZZ���`X�H�e;�WX�J� �[.wJ��2xZz�X� �T} ��&�LW;�W��W��e�.X3rF�<4�܇����*J����*H2���6���J����Y���'Y�Y�� ���W�X@B=;�W�q�?�Vb������X����4s�>b �3q$�B��W���W��ᴂ�x�D��8q3�4�;@���k+�2�D��E&h1̖D��0k��D��4�O5�P��Q���W9'X�����8�N)X\D�@@��WYD��J��P��t�?���W8�?X�h�VE�L���	W�����ᴂ�h�D��8q3�4�;@���k+�2�T�h����W7��Z�h���i���!�TH="U�Zt��-s�;Ӊd�'�W���ەw�5��HH)Z����W���W\����z�e+��Y�~��*�W���W���W���W���Wm(�w�{�h�_ʊ8�WϮ�W�CH���W���W���W�n�WϦ�W�Ҋ��^�W�õ���l=�k��^����,U����RfX�ɐ ��d���<�xS����xܧ>b��1ԯTI�Ґ�1Â����v��H:�l��ߴ��Z�&�w�O�# +F��(�j�J������9oa��3]g��T�*�lyh����dw�����Z̈́�]O�?g�|�{��r��ws��j���8���/��^�t�d�0/Th7<�֦��7��T�]e{��Q�uV�Pt�Z�Wu�L�\b��h�g�c�0`��t�A�B����`���>����Eʧk�q�њ�qʧ��P9T�a6@�5�Ư��;{'}��C[�j��&;�6��ڟ����6\��z������s���_��ق�8z�֢�;1mi�>��s�+A���.�A`���O�c��*I�`�����Ycr$z�� �3��{/���r�A�f����"|l� �h��aoKߧ�P�K���<Ed2��&1B�%�D	�}������x^�[�X�����8���2��z`[��%Z��_�Gm�aGs_�c�x��3��Y��L��
p�j��{���jQ�GA��I�́m��x�9�������F	e!��������6�ox/3��`B1Π�y�a]Ft�#���k��^֯��Uj��#L�������D�K�guZ�}��n����r�P;Л���4u���P37�8,�B�<�JË}Er0.���i�;��ޡ�n4J9�	f\QQ��h]L�T%Z_�̟v:f��m�Y�%.^�6��N�MB�B�$�C�I6=�y��K&���#?���d�+.�i9soW�%�J��,0Ĭ�B�'��N��+�'d��*�4J�)��ʨb\E���B��(>&o���U"�ʧ��OY ��߿��Ҙ��;�מ�{e݃1Qe.�] i����OH�˨�&*i�W��+��p>�Γ�`��v����3�G;S\�Jul�w�PߏCذT���%Y��{T�/#D�n֭�5B���P!֬��Y%R<�X�X�t؀�X��6�<9	����H簭��ג̟�Z�6�,B�u���l��p~ExA�o��8���J�CW�ˊ(߶���4�E�7�?�tpWd�,�Ԣ��]�ݞ���a��jL�|<\�;�_S��������̘�v�hM���ѼEe�!����&�IQ���P+W�#�[u�Bk;��u-��9���O�^�cLm_i��s���sUuل��?1(�Y���
r&[b;�]!���"��#a���6e�Eo&�N�jo��>��L��y5�s]��/���&����4W��T{�˘4���0�۲�TkS�difj�O�j+&������Am�|�&�&�yV���;�3�0<�Zi��UOz��jL����R�U��R7�� 7.`j̪�ɴn �����?�,� �ߙ.�bo6;<!��s��_f���h?�7b]�'0b
�dP�;@���]	����H-��޲Y�MY��ymZ�i�d��dx�����Ӛ�+:�Ъvs®�>2������|�`E�����d��`sy8�25�|?���\�)ܢO>�e�f4X��֘���N2�*ڍ��%""���3��:�"д�[	謩'�&R�R���\VZ�����1�֎�/�Uv��8v�q<^�>����DiE#�/iI�ȉ������E���[�M���< ]�r{���O��Λ���fs �ii��G��̨f3�I#�@Ñ��xB�G�:T}4�S�s�A*����3�FC���x/�`�t!Bu��� ԋ�_:\�8��WSF2 ��eΊDo7��x5��)��N,�Pdƅ��(�wjZ.�hb+B���XOv���]��^an�^/$�Yʇ�\��s`�'K�3�&
�t�s9�/�Q�����f�IU��b���HE�oƲO���s� �H��8<h�nQ�n�I1���Ek�CR�:M8)_�z���$vm%ƭ����l�/:3��U4Z�r�)Īł0��W�^I��	:�����~`�G����^�M��~��Gl�oC|Eɷ�C
W��l�=�Y���βT���j����y1�\l�?��T<h��[F�\�E�`"��T?�������	~���Ͽ��1w�GR�̲��ڼ�/�_����)��,T��5#3r�g���.Z�eA7w&��)��t�Ejy��C����ѧH�4@W�t2����f�"_>կ�ş�QC�c D0�8NjMy����=~�z�?2���1_��hH&<3"g-�����FW�Բ@S6�Dp1�۪�~[Tz�}�ii�@�?9n��W	��"d�h֦,��$�k,�nlwe|	o;����=g�/�ٙ��R�bYNg��-y�P�l��Bo�,��&q>vZ 8+g�ؚ���w������fS��B��˦�WJk��[�j����g|�5�ot*�3d7�K��N]EFo�3�`=+��n�7Z����~�mf�s�E���)�[��� ڗS�IK�T\�|@T�ڌ5u�v��%�!:��zͮ�T4+d��1d~a��ǘ�0r�W����U^��%�9��ρ~,m%^e���	�+x�QU���;��C_���le�<��z
�B	�EX+uKb/��{ө�}�����c�" �� ���5���@b:�Ŗ��d �A��΍/��6�ڨ��]�l0t�ZC$���ƈ�M�p���	�8���̘��*���x�M�2Fz�(���=đ�m��Y��
�{�TM��ӶӖ�źm��芳Z�8!�=X^�l�ӓe�7P�Ԣ��~��BU���[���1�>a�'� ��^,S�{8J	�	m�"���3�VQǉ���%	u��0� �+8*��^g9fA~�P���c/�e���8:(rS�n�^}�ㆢx� '@��@�7���m�L�k�x&j��cE�-|�^�=��q���3���`�P�4@S��$�˥$r�#w,�ĵ�O
�|s8�	�x�r�q��S���v䂴f����m�q� ��' j����c�C����d���x1� ��B�.�E�^��)j��`wS�Dw\dLG�S�6�
!Wf�u����q���شt�[m�#��0&��õ�|���8�+Ρ\w����j`Z�q5�����- JS/�͏6�� �HT�ⷕ=B��1�j\e�t>X�@U��n,��t��=�l�<�Kv�	�m���Qu����g��Oy���>�_7��S	��]˰V����<����FΎ,C�]7��X���)�ޭ�[j�`�}}Z��9�	l����
���&1��N��:�
�y5���g���ie�44�|�~릐q[��3lxCk���B�d0�J�WN ;�m0=Y�^`��N�<,ݪm����3Iv}�������T��~ii�� e���l����@�%?���u8��bΘp�~���_����E���T���A�������t��w}��?;�r�p:��YF�*L�ݲO�(>���J��rΓ��^י?m�s� ���]v�d����?ѕ��ْ�"z�����W�",���֟-H�:�,����$����}M��ի�^���Y�������)m^a����p������9;�O��l(�{V�~:�B��u-M@��=���*��mk��!e�����A���c���ƚMr�ݢq2���9��p���Я�<��ڙ�3ʝ��Z��Yu�#���"LeB�����2��k���/�к�1n.���)b��t9�E�r��(�F�I���Ͷ2�&�*�K�]��V�*m[K����������Ķ���$���J�mJd����vr�Ю-3��Q"!�4�?6�YY�f(xN'O�/+b����7�%C�9���X�Ka��7�����2�ц?�Z �B�m������{N��ʢ%�v��{����u�3Z�~���'����H=ȥD�Sܼ�eF�ɠ�7Ir��lҕ�o��:�@��v���9�����)y'�F�0r,�:u�6���`�˝{ZP��	�CJ@�B��y��d�����a��_+-�(��V spo~�x���T��~��6�pE�8��13�{)78�l�S�k�s�\���
���r�D��8Z9[�T���9�5�R@�z KG�I?��6B����`���SДWIj�e�J���`'(6j%�q����'�1̣B�Ĳ>;��$Z���=>��9~�<�����OmM6W�߅Sq�>�t1�~�z���.g�-F��_gǤ��� P5� �.hwR5��[-��*Q�tpO{�9,V�V��=:��E\T���$8⊨'�a|�:m��QJ[�^!w���e<LJC��_��ǋ�)fP��i��pΒ��RU��
5r>���I�ɓ�"��a ��-$��B���K�~�6n��qnt�!��h	��?���mKI\�����}M
�^2L����J�u6֩F7o�]��2��{���ce�R���j���bL�� CQ�w76��DV��&N_ϔ8�9��'�p_ia�I���ؒ	�5��F�u+l��MW�I���1e���~��&�m�s(|Z�)r�s�H��j%a�{��)G�$ʃF�h�0��ڐ�Jf
�q���FM�a�F��")e���7r��P+�!�b�	(F	��E�����kݛm,�;��w�������d�y��e߲PBA�+�QRP0�Y�`�.|n؏k�3��(��ߖ��_X_+k��:�`0�{z9����7x�a0C"!����`n�����s���n#����L�q_�u�&��\$��$bΡ�p�sN�`���z )�S$���eF��3)΅�B7�+ڜ*)J�Jy�~�-H^O� w]�@�n�gs��_� �>���B�T�@�%hQ��w|`���*r���	⨀[�E�5�&�%q�vIo�_|ק�sB��Q�0#�*�1G{�T�u_���b�
�s�	2�A����u;��s��*N�F�����k�:� S�r.�)ڑ��6�fC���Ey���>�F�ղ���L�J�4���Tb�p���E�F��vr��yS�DP�nB��&��r@mC���L"6� �D����іD��wp��MMY��tʵ���"�\yY��\����R�pʠޙ��Q�Ńx�߉o;W���QH�D�J���sF&��}��i<�N����`?�[�r'�����Ox�����."�Z����z0<��c@18.W�8Y��zZ5������+ɱ3ή{�
�:�n��G*W�s����CU�.���Hd��$�c���b�ʚ�s����&qvk쥟�CEKZ�ϲ
b(���WA��U�<��믗��,k�]��K=9��*�.�^Ƥ�d�(}@L��Hr Ƒ3ir�)�vؔ��0�n��[,�o�R;��N,ǹCQv��U��ӡ ��~���~�<��0'���7d]��ڞ+hx`�ѹT{6x�&v&Dps��	\���q�6��-%f7��T���(}k�k��Pa�̩daI�>K:��ZI�$ܹ���VW����30o�˚l%�sB���L:f�����~���j���
O&=9IR��{�Ib&�7�ص��T[	0u�� (k>F��qH���Ȳr�J��|�o���2��e�b��l���P��ڢ����;�BU��ʉ�J�^�g���aW	!JQ� ��>򐆟J&\a!�HA��d7K�%U��&BhQ����x=�ַ����i0<���z�+���W�<��gC�sT����M ���6.y5�f���."�jE�=A���O	�-sp��>�j��(����?�J �~���i}M�8.iS��ZhI�)��\H�@Dב\&_ �� �L;T��Qf�j��I���.j8�q���3��k�dKԷg�6���؉ÿ�`P�D��q�Q������(R#٦]����P���0��(�����;{�����+�ݢP��W2����Y�y��P�[=3#x^��cY��ծj�F��ӗ�����o���〚}��/+ɦ�܆o|#s��6��c�8|��"4�@Y4���Ϟf�V�H��.��55Կ�7��R��(�S֗"���!���a��Yì��FYY#A�=�,~�t�s��ws6�j�����[տ���y���\B������.����@��Ptr���ǔm��7������D�`�
8<4�$�8�׵an�;���{{��U.uW�]���t?�S%�Y���/p ��y�u�m��8��/�Rp_#E�MP��+U�5:�8�&�g��χ�X�>���dBL�
*�/]�.�+�G}/���������G�����h$���������=,1�Q�����fz9�Yߥ���qy���[t��W4�.a��l]�Z��@q��4 iۧ��(!��vB��a�Qk<XW֭N�ن0�P�gazeI�'�-�$�civ�ıA�~K��]U�4���<�VN��/��#��_w��k��熍�۵ݵ�7��:�VsQFH�TaCg����wuNh�ۅ�H�su��T�^��QDB����-ݑ���ŮA�g��ƕ!�AC���p/���y�Fl�{L^�<~Ō5�u���/ϥ���<8ت,���)�?wZ���]flz����8�"��}��J���Dv��Y�vû�u��&s6d��R
���UG+_���ij_kV1hmI�5�EW���- ���jY��35��.s�d��`>��tR��è"F��_�[jW܁xuJ[�m*慞�ϋ�L�W�a��nw�o��`s4\a�����PEl��/�.���T{�5<����c#��b�s+Μ�j�����˩�ay]� �Q-.5���J�z���#<.q��M銅�d��y�pY�9F���/����������L�Ǳ��\�L��N7�&[���� ���*B}��!<9bN�� Q2����s�GΗ�g���P���gpDHs���3oĬ��Dy3�t�c��~5���f��Y�*��$"[J��t	+s>�Y�zI��9:��a?͢�a�S+x_-H��HNd>r��}�j_~��MKJА}Vă����%kU+�?e�5tMF����$M5�?}m�	�.bi#�T���r��cZS?���j>��Hi��W4`�W�l��y k&Q��+9�^ߓJ�ؘ��2v!�<��{4T�B_�5����w1(|�%�n�ޯ8���)�zat�)����w4����	��=NW��� ������/��:6IU���)������@ä�:�=u+���pmqǂ��u 6��[P�ʐ9	����k�o��>Ҫ�XTk��G��Yl���և�#Qq���@���������"N1�"�nF��%�ԃ�?���S�����'+Ue._�A�i]1F���Ok}���~����Mk��5���Rs�Oؗrt�y�(�'� �l�Ou��$ОjA�!3�u�\�:���~�F_l��k��z�E�ü~m)$=����-\��;,&-�x����:�P��x��i����_�DZxHI�/R��u8�1,T���bY��������}Y<l�K�b���=�e;�6����fx���z�Z�M�x(fg����v���`��[=b�q5��b�� 2P^���ʃ#C���M �;�U�9��H�Z�������#̭&;
�@����临~��k�&��CÍ���)c��V��ʱv��!��F�;0����O�|��ͅ)��t���o���l���z�	�䥋��j���i���y>��!$GjWܞM�)��e����[��u�0��XSO`P�F�Y�(\�/@�q���J 9�x�T��ZJ���F�'S�(��HjR6Tn�ն���i��i�a���Ȋ���vleB�KE z��A��&�h}��$�`�^Fę���,����2D��௵���&O.by�8R!�([�V1pA���ca�$!m��똝bi�	Tƨ���Rw�3��6�,�lnS���ciYi ��dM"���{:�ZV ~l��^(��&*V�:�)�c��r)�I�l�]����a��*�S�ϸy�K-?�}Q�Q��6#�Ѝ|i%9Oy�$��3Li��KqW�?��C�0�aI+郂r�?�W������� B��Sb�#�K�@��ʱecAm~ 	'T=}����Փ���윰?hJ�0%{�#��b�'�?�"|�U[�(��{����xut�H�u��gq����bH��N��%�.�L�#�8bi)�o�r ��;aERx7��D�Q�d.�N	2]�,�����äO5m�����m�ZLw����_����ه�u���5!����՗��|�U�d�ls].�����hF�����k]W~���"�$�)��[<�_	�}�-&r�K���u�V|��<�gY�޿H@�z�v�J�x8�P��̫+4߬'�����!LJ�'���uK4��lN�W�&g�-��js'ɦ��35��x�R�=p�x
�3(���X�YݤA?ԉ�x<�`����M4e^�h�T�WIE�d����+Y�M��c�̜e��贱���,�Ij�A��gPF?d�"�	Ct�>�ߪ $�۫��ae�3�	�)����=*\�Q����o�2�&�Q��n�%��1G���٣#$���uҁh#���0De��u��4��.`�5�̋�&�1�ˌ��.�@&IQa�Q��>��#i$��{�N����Y��u��?������{Ms^����ˍ�����ݠ��G�F;���OF����C�������w9@��������Ǎ6�<o2~��m���-�S��y�rM'��5�H�[3�6.e�M>�-o���P�g`x7e��~o[C��an����ǯ�~W8[{3�	�y���0�+;D⿓�m�����*׏N���!�d�	\���H�ص��F*lo@�n��{�.�m�d��GO�<�x�1��O���[����z ��K�����5N��)9���͗�|!s������ߡ��5`SP-7��T-����L�4���@�ʼ$��$T;��H(�=�؝�b�>��0���ֈ�)�SzF�LH��������M=l.G�����i
��^>2��|F3��͞JfHW9�+�Tx1	���.�-�����Í�Ɉ��+\��)�2�rE�ҿ���q���2�%c�3X!�S,P�d�S����V)�� �=Ylt�Sv�6RľAG����뢶K����V�1�-a��tO�K�O6\4:Ǭ��Ϳ�H����G�f��6�~��0,.70�G�}1�/E�?���ܺ&�T��$[��.���)bo^Ӥ��(�����U��xL����w�"�`��R\����Z�Ho����w�x�9���r^�n���Tl�BBa>Z�ԧVT^D٢T����h�D�9�>��qKh��������T���*��������^�3,!���!U�X�l���C\J(�ڣ|�7��J������
K�͈��֝��Q�gS�fWܨ���{3�<$u�R3��U�#qق�̕n`������������R�>��?�����g�@���q��˧3�D(g��]ce.�LrB�N�$��Y��v�[,0*���o־|m���w5�dL���ia�}=�q�w���G�/1�[ְ��ߝ�m~G����d���S�Cf�,�����k�c�lŶ��NR1m�h���z� �U��1�n��s��YH��[_�;8���B�\�END���A��ћ�;-J)6_�ҷ#%`��My*��d�z�yv*[�֧[_\��S@(qj����(I#n����C9.�k�~F�TN_\5��/h7eF_7�-iuͺ�:m.�f��U2s$���J�������6����5�ax�(�8��⋬p#�?�&����$�U����Z��M!EJ��h����PS&e�N	�[B��2^�l��րJV�w�$�ᕂ�)q&��ҙ4f�F�(,A��_<�Vʯ��(
�J�*�4�^��D��l�|���G� 	�~N��.M�R��{XS�1��4����T�ڐ��0c.�9rP�b�pi۔�#e�ݹ�`������y�5Sl<x�m��}|���X2%8L��Vi�߷�i�-r/�u��X��k�#3!�ic�fƐ'+��ߛ�����7���"{v24l��\�h1'T��@�5���!��۠	 .0���~2^x#깆پ>���U�ˣq�Fۅ�L��N�$=�2��!jg�g+��_g�7��U�F�tx$�;��V��;�-֎���ĮrE���M,ڻ�Tj_O	w~??�*}F.���<�F��D���]��!��G��������}EN���r�DY�eߺ�b�QC -��R%a;��h�"�"��}[�=����A�q.p|���_�
8P�C�?�V�{�đ <��:ν;>��[h��K�V��B�y��`Q�]B��,[S��|;��!�Ff�� ��7f�j�֊x��^�j^YDk�	��d@r�i�hEv�.Q�#�*a�����ZE���e�Z'1�^�^x�u2|y?�M��&쟏�s�am�(F���ƉrA�U� ���̕=�ەC��*�H������;��l�� 
,�U��ھ�P���o�L�>�6���|��H�v���rn�:��S|e�x���DԄ�����aё�;3>���=L��(z&cB�BZ`ќ�Y�����z�<p�����F�W�w�i�<<M���Y@�9k�MA'��o��6
~|\��I�ĬDB+��Qs;&�k����Ƶ8ĠC���ؼ�d���ʝ���n�N	�[��q� ;�t ��@�aqjb�m���3lp�T�N�B�p3L��Y=�|7 9�y:Qs{8[��gFe'w��|S}{�\g�ߙ:�E9�>�ʹ����t� ��J�������yR�rB`Cl���fղw��=��Q�5N9�՜�P����8���텎��%��E."9z�������l,�X?��#�\&�σ@GN�͊{���~N�1�d�H^�"�g�V�C��q���v�׏���xF_<��#�w~�ʕ�,FY�k`i�C����^G���C�E�Tq�VKY��1��R�k�C��֭��IC����v��"�'9�J+��"-�y�,��/Jי� �
x߾t3mH�N�e��Ø鰂MD���(��<���WH�.�Ϙ����r_L/ᕽx�-�M60d�j��I�O������F�b���@������K��n+�(H�3��.�� �I/�O��7;��a���[��v5�șo8N�%�*�`�S$��m�V<�	&5���qA�/�F3Q��]� Hz�R��*P�պ#��~�6>�L��&6��8�gQ�i����X�j;�&}B�A��W^�����N��.��j����Z�؟���k�:��3��xn���V��~�?�?`ʻ�b\h�F|W����wN
�������_P������'�&��UYX+l=�W����o�/T֛s} ���ƛh3L�#� 0{B �_֍�}��<��jH�A�eIu��Br��ښÂ���?)��&Ӣ�Ƕ�`5mK\=�镝��c�ϣ0p����q��9b<�0�V��S&�~�ܿ�y��������"����p	#s�43|�h��y����+�/�Ҥ����0���������1�!�Ivś�7��3�_��j��cquR#��w[�>���Z���.�萧�I ����A(�r�/�2����6�}�P,����f�`�e�Ԩ�H�7�-�H�ߠ��#�op������v�D �����;�^-�G��I�AS�4��{}�i� ���!%���Aڃ�f�'5Z�r{%��Z�l�,@C��3+�J��$�(�(Ղ��E�w�o��z�D�PR��R�u�x��^z�=P@���cK�Z�JQ�K�|"�&���KI��C{�4rP!zK����P�ԞRA͑7N]P���Z7Qس�1$ ��=J:�ŽV=���P�(��W#���\P������])\�d���p�Xvb϶�� 8��vƉ��u���JH���sbP���h��
�ːb!W���H��?\;z�n�(�i[0���a�����+�Л.�m�Uj�S��,�@�.?k��,0P� �/�#�SP��t��̯SbU~[7�H�E���K0�g���W�O����G��	�d��^�J� h&��65�4��,�����%��j��"�n��y�����8�0�@��r����էr;�2p 
�a�gD��`Q"��{b� ���&�3�G�5Z���>��ou�Ғ���\�����>N]���I{D�W�`^���#BRr��=��.�������H���J��59VvERD��A�j�9Ϯ�r�p�@1J�5!�Z���O�M����2��M�L3�%U**B�H��i�>.���Q��M�S�Z�hB������Sv�j�sk���q�c� \X0�G��r����\L�u�'�_6��	��^뛴�̥�k+E$	.X*a����~ B�
�
����ۦ����V?��m�GA��bF�ԩ>[.�idgxQ*�u����S_��7�C�טvUe����&{N���?�׭{���5���6������5da�(�	ts��x]|%X�JUg�F�����C����+�b���+���Rh�o]�u���/��˻	*�F�ΈU��ڷK�j��U�A�b!�!Q��ug��e� �T�N>̟Ш�7W�_� �;���2n㤍�#�?� ��:��⺊i4'7��������T?)w~�ǂ}��N����/�D;'�|������`�bW)���A��G�ٍ(p��O�.@����Z`�R'�PTG�� ��y�*e\]�u���E�����ҝK�ҝx[X��9`I$5M¨�^{n����[Qb t�d��L�ū�w����A_6�+�K��r�ڟ0�{��ob�H�S����
ԅ���z�[��X��`k�zg��66���@ %R���|�!:9{��B�9�|����'��	�5[a��P��S���&8�V��Df]��A��`�>H�l3�PUM�f��HA^30E4���H.��H���WC@�Y)�l����5ݭwv� �w��x��N�}RxD�C����5덣� �~���sz�wq�|l`p9^S�K'^0?OF�x	�(P���V%���*�.���S�B!O������/|y\ģ�)�i��l	�@��s��H�̲�]%R+	rySv鳖A���VH�U�>�k�pe�$�?m�7䞂崱d�A�eHg�'F�c3^�y�QE�v�Ureۀ�W�bWq&���>Pܫ��m�zI�W����D��L>� �Ѝ�C�T�O��Xw�c/U�<�b&��8N�s��������8S����Z�m��B� o�p�� �>P���T��>�/�R��aαd��}r�ߌ��(1���p�e
�T6�Z�^��NӻJ��t:�4�t�� �N���~Ts�B&��#hx����}�|�oQ����9�e����	a�����
�)B�)�0oZ^�����huz9��(�����,V42���j,�+�zg�(?=�dՙU�#	
)�S��s1�v���ۥs��^���n/s�<�Ԥ4=s��*~����5�՛���v��\>cA9 <���j"AuI ��ǔ�hS�[&���3��W �wp��JA�O��&��O��frj�ݹ2z���2
{��(���������Ed�����Ѥ,r��G��2
��3��S��vG-�|T��dl1t>*�a`�cyr�}���,���~Y��ZQ��t���f 4�bT#!�Y���=��{3}� ��m��o�	y�H$,�zo���Ϊ!�@4�����ZV��[OnƠ4�@GĪd�JC�-�lp�o� �eQ�U~�+�_D�9�bL��}l�a��:JxM���5:�`Ǻ�E����E���_� I���i�r�X�'�#6�L���T�rS�ID���N��,+�=�kʦy#��x^R_����S�S+$U �\�kgr�:�q@R���T
o�֭�p�इ8{u���"UH9��W���o�p��y؊��Q$q^d��Rr.�Kj~��ɀ�k	�����W���9�O�ߜ���
_mZ�:�ݥ� ��I^����r��Nn�%g8}�L�2�"/��r��a{�c��q^�8�]]Ś��_:�z  �S8���_�&��Z:�j�u���0S�vVj�=�20�q�zގ��QSi��	hNK_IH���9���Ѵ�M���z���q%��O:$3Q9����0��r����_��+���İ������������>�Һ%�E�~� �@�-�{M�>f?�d��ｱgt��P'!��(�,V�w�"%�i5�A�2B���	����;��:z�ьZ2��Ŭ�>�x>�tm=�ߪ��h��%|8�.����N+�Ş�Y�E|!���#��ZMɑG�}CS2�t����l>~`�<w-t#i^k.Ѣ�=,*���~+C��6u�>��4��.GT�.Y�O���}���hy׸����^�Uf��披�w\�)m\d��Y5Q5������t,�܁.F�H6)��w�~}r>�Bz�s8d��l��b�kKء:��B�;)s��� 6�j�?�K�W��3���@eea��(�6�Ǖ�N ����F���ɀx$)�&̏NV笔	���"���	3f���ҍ���Q���"���h��H��g���XV�H��N�ie=�� ��G�;��#�����`���Z߸�����Ǒ��2s�c_hO�O��]{~�`*��;���&��t�����)�$�5��Crs~[֫�䣄��`P[���l�?<�%*.Ѩ� �Q
VjAu)��ᑑ{��s�y��⦦��]_�8	��Ů��P���q$���i��b�'��M��尻�e_};rӌ��Y�q���H�)�PHf����5hO�$jk'ny�~0�p5 �j����6˥��ga�
� ]��w��;��,pm�] 7�<2����f̥��5+���Y ���e��b�Ӆ����_�%��r���jw��]�����=�m�u׫��Zi�
Iɿ�?����"����^��%D0�h�����s���V�1�Nh���؄M����Tz�K�D�����+���] �[�`����� �p? v�\<���vC?B��|��y)=2��H���#\����q���e��S�6�-���,��Y�,l	�E�:�p
��\��r�(��i}�}Q����;�	�݈Y	=� �ʫc%2��1��z�ʼLx�#P�S��]�L�p�t�am�ڼ�d���KK}���Ө��pI�~�0�:}���s���VONUq�V���;�:~�Q� ��)�i�x�T�/1��{�"�$/agH}Y=���bWpɈ�ѻ΋�u�Q[���92�k��ǥ�=�
�7 ;,G�R�~S���&T��0��0��6�bAv���k��Z��淯XX��ND/lg���#�����k�U�G v�qE8h�)��Z^�/�TM����gI����m[�+���d襉���m#ˋ�48L5x��`�������<�f:w�8�Đ�+%�t��bs&ob7�y�0Q��,��;���w������8~���|X�υ?(��Ƅ�_^�.���MJw��Q�ҹ�颤Յ�� ـ����-�+�N�8q7{+&m�J�,�b����*�S��H��>�B��H�Q�sĦ��[�0Ǳ(Sq����ӵq�fq�H|E���ު��o�b��,]�A|2�_���ՙ����X�N�[
�@D�o{�T�+�>J�Z	:�IW��a��xj|c>�=+������!�ׅ�b|s��wK=;g隲��?�F��y}n(�c�*x<�:��5�b��ޑ��8�B ����R��u�x,g�l2�~W��'Ƥ��7u�ΐ�Zҭ�j����;t�KL��R�Ŧ���dyTȒ6}�r��
��/^fD0�q[q�������H���qM��Q(��G3��v��(Wv�:���h}�EJA>H5
��ꩥ�3�]�t�5��э>�����uA�B���-�9zA��#F���h�� �̐�o���1�-��7����J��um�����\���	�Ƴ�^�I8F�~�	BkF���s8�H=�4u!iK��
U<��f�:$���'��ܽK��Yq��Gԟ���y\�j���#rt�d�Y�%��4��\�x<�5Wۇn���r�8<z��h�=�~8��]�]�7���@��	��r���!)Z�������B�m�^E�.��Z�|�U��0��M��#c���[1�O(g�<��c:�+3�dE�lW�{afYx��ӕ�9)3��/rq"�:h[����*'c.c���ƣ. �I���u�5C_n�RP��G�QH���J�M�'�9�^ӳ�z���T�q+�~��Y�����n�xk���IͿ8���\�i�߭�~n�F^�Ua�P�G2a�Ѯ=W�r?�yR9����_n�3��Ez���_[�a��%�M6{���3 ��J�|/�.���=o���M�|�`[%	�YJ\�vv�b��)��Cvݦ�P>Nd�x�G��H�bHC�c��Q�IYHi�ƽ��G�Ξ����:	Fuҷ�4�'��0��_X�>���g*���d�1�1\$��o'1_JŚ-Dگ
��؄�	��q�.O��/p ��B�LL'��F��e.s�����7N�_W��\����{�����v�����5Db$�瀪�ɇ���!B\��g#}z���l�UJiuv��&n���-�>�S���Y4��l�G������ׂ���>TN�%[ळ�Yzs>x3�DX�#��U
�d!5��]��~}lHZ+RA{r��f)�=ܺJ�xo����azFQ�*��a]�Eq�Jo��zϨy�s�\��n�=OU��ŭt����:�����Ýc'�����ݑ߾s��ii)�}��8VK۟yMPI�$�SR��v3Ulb�hÍ�P����vcY��.���Y%�s��V�[ q����Cԅ`8�2X�*��DH����YQۋh$'��6����&2�}˖��#6���3��!�*�*0#Y�-s1DƓ�w�$��?1�=$v���[0Y�X�%��چ��YI���Cstk�;�K��'�2��H�����h�X�_<2=���X�ՙ,�ZG��/,18�|y0�8�%:�-)�!�<��e�g�狗$?0�~�:���{=���O��Ö�/^��
e��*��A����<Ў/��l��2�R)I`	.Xdor�+��z2�^�CrvR:���� Լ��̸�u���k.�@f/�M���4O�Z��YQ�^fwE�9��О�]Sq�E5�a����ziT6��K(}���=�" �ۍr
�3
/S\��W\��72"����d�	&�W��^�U���^稙q�b՟��!�ǰ!Zϫ��x-�$�((ߝ̾����t������9.��k�%dOJҚ;5/� ���<�sc����`���J�9yQJ�S���!��D���qF�R�,��=@��4�f��]Mo0��m�n�ё�D���ײ�NV�&��:7�U�%����A�xK��cK�$��ٱP;���sHg��12���� ��͉�ܶ��ye�|�~b����@�.4xe*�g���r�-��#{t�T�� �C�\���9��� � �´�pC��o	����Z�"��k�S�w.=���g+j&F����q���u�A��bK��i}#Y��<�҄5UY�S���<�N0Z�G��`k{JjJ��ȸK��G
�;��j�83p����'�T�ʂg�g�����M��H\Ë�B@`��Ej�0��~=�C�����_\Y�s���NH� u�z�W*����|��@T�5�ܵ�	��Z�A�{�t�O���.	-�u�W�E�����q�� |ZU��ȏe�1/�P_wmk���S&��`�=���g#�[�9C� �i/�KA�b�����C-�?�d�2��`T�"���2�s��`x��f���OӮ��xIm)ʜ��j��8�J�γ������B�L�]����_����-L_�&�9���Z|�.���T?�B��a���t��0��N%fh{|��0\��P����-�ڊ��Q���K��6q�p�ߟS����j'U��ߖ��s@�?��֖6�HY�ܩ�K8{�P��p$�T\�X�x�BMG!�u�ҏWy�&��e(?Gº� ������-:_���U@�m�%d0#K�p��h��at��ޥ�q+.��6��쓇����mYtB���v���dhp| �$�R�T:�����G�i���+��2
n����3K/���#�<�N�nc���)���}��p:�

p7�]�ގV����*ri�nw�fm#�[W�s���G��g�N��x���t���bĜ<��lzb��VO㋅6����&��0埋ۑ]o��?.��V1W�EU&h�p8�Q#�R���|�,�CC+�:��w�wKqo>;�h�ķ3Gb6�2���6�n�=�o��R�=W���gˊ��w�K\%���Y@X`��Kw��G��VhM6I8;ь��Πy�+iΰ�P��rp����'CfS�& �a N�Vyv�cd����,>��qPQP�F�Sk����gi�w�6�7RQtf�^�亖�,@�ܺB�1W�JpR�t�,�F?��&��	�;�؈�H���H�EW5���+���1�7��E̋���AyJh�}�X�W]o�s���6k����PH2�w�V�)>�~:��L6x+���˟�?c�LZ�o�
NLrF���@�WS
�=�w�,�d��������w�ț��U;� �TL�B�$Q��j,�g�\�/�"8O�k��8Wg�x�MF�������$�^S��Tɭ(tLʘ{��+�����V3�b��U�/�_��Mh�ZӶY3Nܨ1�L��<�}=���������L$�{Sy�&��7������3�I2��a��(%0a���-�p C�
Jrӆ��1���#H�#�&��Z�� =��j��'���S���f�ɵ�v���'��C�����9���OnM7���d �uY�Yn!���X�% �b�B��	أ !L����R��!R��;.��:ذ
n�[����a����i˞�!ѝb4����l(AU��g%ކ���	9EI&�Ք��J֔���׮D���}Z�Գ�����x����&l< ��ya��L��1oȴ7㕸b�f���I�$ɒ*;V�{LK� ��Ο�t��Ju5����4lGp��
�P�ٺ�������׷�V�-��Fr��{l��ó�N�1)��*��
Z��GN��c�{؜����qr�qF�i��
�Kߑ���Y���Vaw�M��2`q�o�}�1u�F�
 0u����j����A@��������cr_

���֞igE|9e/�j������]ؿ�U}[;�����S�J��9Y�~܆�g<�"��i��@
(!�$��i3f�Mmj����2v\ {�=�h<~lE��a��_�}��g��������^a=3j
�Qr]3^10���\g��,���� ���yh�eRJ��8>B�G#����\�w����/ٚ9�q�+�!�h7"�3�����G�n)'�l|�3c�׆pm)%:д��cX�n��)U%p��X�v�9�����4}��
?� v����! ��E�ђrL�[prj�~g֝x��3�r�@��,������,)V��2��C�T�f���k<�>=Em"x����p�4	M������ˆ낂���9�P�zs���|�?�^G�D]&)�B@F�J 1"�N����;����C����mH���1��V���Љe��� t��5�A�a��A�QX&"���B?���b�sVg̛��\��9���xC�  :�6q����� ��ӟ᥾�<����2��W�VHP��mۭ����{�����C��nN�r����	��(�~)y���%��,)׃0���u۬^"���͗�E(�G[�#���]�k���C;%���E�b7��▷Iv��6 �-�.���W���E{�暟�̀Dd�>� (�!�?H �U?~`˨n�iy*Ա�d�����Tr#��w$�����#Od+Ht�z�`֗�X���bS2�݀�M�z��k \'��!6+S��F�:<M�S_�{{�aCT/�Yߕ!��f/�i������͎;��_G\�y���=�-�lp�E���������
��?d����ޜc�<�rC�@I�Jc	��]�����	E	+Qorrcׁ��t���߷�9Q��u(^�GP�Z-�n��M`�u�wj��F\��htc�?�F�Es�|V%�D�A��(�mP�}��i�d#ZD�D����HV���b�"�V�5�zR��L�%��ア�A;>�|���J><˵V6�\�A�tw΀���2���5��9 TQ�����In"R&���&k0��៾7z`����n���Z���-r�Z������u`����!�%f�/[�OZm �'`��|����5b�a��P6	���&�_���Z�����:9=>����f����
2�אs�6f��b_a��VJ���ΰ�LypRo`jTK�}q
x%���HM1ύ��+75��K}ȘF|�׈��b���7�i�X&�5Y���Qy�1���4
�/�gM�,q��ü�JP+@�æ�������p�w�"�&a�Sȴ0�@&�l�a����a�	MS�^��뼳��x��ʯ¸��{��Oիt�'@4�U隸Pi益A�-t)��rQ��b^a�5��g\��?~���7�y��[�a�y�R��*!�S;D�:Q>Ʀ�zd�	X��1^�
�R"D��#z(�Ј,b����Tt&��6��7 �'�.ھ���g�sh�?h�Y�*k
H��Y�o�T+�����8�.�Gf>m����t�<�4�׭�r�z�*В�4�����+�e�κ�E�n֮m��\<��Cc�ɛ�`������{�o��(�ɕ�",s�\а]��.��p�Jum�R[?-�j\V��CcbB 0����]�"n��ے�O����|����,�̼c��,̚|����햯/X���)�{½��yc6\kT����E/~1�,R��l��HÂ��B�t�0N�p���D�{��A$L���r(j���`r4�vje4 	��6�(2G�Y\�;О�`�49t lN�ޭ�z\�g�%t��Cv�ŬI��I�h�z���8��������퀰������B���m��${�1�W�O�P����4�칬�_'�`�|������$O���k��|�s7�q�;�M��!��Y�W��'��'����o��u�?�N��.+����&������ަ�0�A�6�<��[Q���
3����0���]��u�
��g��Ӥ����tTe*�L������!���\� h���A����[e[�</ �7�[�;��k r@�.&��;z�έ�A�#��ě�u�Ǵ�������@$=�U��t�ɰ�P� s�?l�I�z��xp�t�]��6�����V���0N%$�ָ9؇~9�C��8am|R�����pyF|�.��`p:�*S�@��Ɍ�o��[��c������ �� �������GV���v	^��M\�C�[:`�.�"X�G$w<�Ώ�0.M���u�8��U7ڇ^��N��_)���{����Sŉ~`i䳥�lNf��T��pmY��J���Fdk�wzA;��>��`���r
Zɮ�`��ʀ��{��)0ݞ��Qq!T�wQ[�~E2�]��V��<)-��*]Q�fK�`�נ
��	��Z}�wqI �oS� �=��б��!������D囕(B��GS�a6���b��d$Zg=�[+������# ��@4��}�`���|G��Gs��:�m؄�Q����ʄ �>Q���L	���|ȗ��#���2h��Ӭ��'��f��X::W���T6Lf��yi{�=�Wn��� d�e�y��J�k}�_�&7�qs�2[;���sD�v�T�/?g�m[�L��I��>�o�IB_�%�����H��{9U�t�hHj�t7��n��F��}ƬE[���V�(��c�e�q�K����3|k������`��j�&������l�n�PG1LqO}�l_�w�!�|k�v�����y�i�
F�G���nM���U7� �.jF�27|}'���'�j%_���E��y��d��G~.�ΘEʠ��՘\�V	��?3�e��.�&/d}]��;KIA��^<�~�	���Q��B��3O�p�Tj�b�\��M�T*�5v�8ӓ�o����؆8߮�LxG��~���~���la�}�8m��� ��3��Pa�N�%XO�ٺ$�U�H����~H��s�Q~n�0��'gCS�i�f~��_��0�Ub%��� ���Yh���ۚL�s��X�ޚ�n%�k�q���Wï�OQpA�Q~���ʹv5K��YW{��z6>����~נ�RX�|����|�l��X�#B�]��O�N˩���	+��7��I��x�4aE�Rꞓ���L�BsB�F��oQfowQ�$;w��ԃ���8y^9��=�!w�Oʹ'���B���g#2	�ɫR���FȞqE)���\B��z��� �3�\�Nsn����B�!IU�t��-���8=����'P�"���Y���D�-�I6F,o�S"�il&�>^T:�58|�%&�1yW��K�E�#�5�tc�i���-�â�^{�'��Z[@� /h�P/�#�݉m\�6��
͵ʹ���^��W]���.�kF�Z�.c���k�2M�y&�&z�D��ϟ�r;n1Snl3z{B?���pX3و<���La�p�����H�j��C$>}�͹KRZ��Z AD��y��>���`ߤ�E�S�@��g���˯&т��������/u寝���hD�r��+P��Hb���(��фVw��-;�K[mOGO��'&�"K�Ϗ6;1��;�Eڵq ״%���[�-e�F��+�R}�&K�f3�e���[��8ي��1�B�TϨs<x���_
5���Z0B��輶�).�a�R��5U�5���t�ƣ���8y�!��e#a��zM�-]�N��ក�`~E�����5���_�����M9eYf��i�ܡ=,���I���4��x��.y��|X����d�m��(=��/��N?��U�5�e�3�B�[�Ţ�4������^��ݣoS��*CN#��]�N�R�ڝ�x-!.�I��L;�L%-�@�}�M�~ A2v��8����B8dD��b!��4~��t+��RL$J��L�N>�K�g��:��1�Jx꽱�T�c@K+��1�	Hz��}� �V���-�W�ثA?��f����â����{�YD��*�.8
0�e��74��bZ�EY��Q8��������f�A?���[�Xz��[��a����Fd"z{���/��2=�x�Y\��J����
��]8.7]����ʶ�C4��Sq��f�'�.���K�J�Оusi����9�C�L73�i�@g�e���v�Qa�^�<�q�����X�6N�Y3�֦^�I�����m'Y�`��)T��E�[G>�^;��<��I����I��L�X�+��x,�Ƙ�O^��[ĺ
��R��y&������I� ���$��3��? ����?Γ4�
G�1�S`��Ҕ�	h�Zr��8{sq�E��!ū��q-��0k"�ɡ�Z���tR�#@?�Q�Ȁ ���#�g{��aCpr�r�k\��Hj5�̚�*3��K�xI(ʛQ$�Pmkni�d���#D`YR�
b#���27<u\�SR�j��ҥ�[}0�"�����uHΑ+��ӡx�K���ȨD�Rw�a��(���ʨ��F#jC�����
�R*�:�o��t.��t��q���?�{�ׄ��4��4֍�3���a��I-�,�(���rL����l{��A��]�s@�0�=�1�A��E�c�e�B�0�P	!�f݁�i��侊��[䲹��Y��A�Q�7�YR�H2r�`���y�N�n�=*Nv;�������v�=�(l�V7�P��ų���K��ʱ	G��n	k0�oL������g�)�F���?�ͫ8�d�{I�J��1��� ��=�^�h<���J�Te*+n�]x��>��S'��)��՞Q��%{[t3���'�*A�䈰A�D'���9w�j�rͩ������ ��ܩ�vZ�|mT�8�(��j{^�!	�����g�����4q�0i'Z�Q���]�NX^X�.����9[V�����oH�|P��4mgh������D1��N��p �]J���q�Q��g�wҲ�D�g)0{.��N���vz���m���I����ՙ1���*����J�۰vY���]t�'Ӹ�/��<EށDXU6w���]����ktғk��2P��{��黠��Wbqs���D��;B�����Q.Oon���U�K��B��`0�ɞ���2�P�����Y��Bbp�5Ů�A�$�����zi�U��Gm�E��|fZC
x���!p���ܔ�� �]y�'X�=m�����Wg���UO�<����#��2�Mo��.,�������^�ZCZ6`P���b!��<�_)'W��U2a����M"�V�T�Gd!7yS�q�ӆJ�|����!�e� �%<�{)6+�/�T����> ��PI&��  �PU	��=ʶ��<��?D��q�M�-)���cP�u
{u�I���p��ơ�����9�/ni�c�;��o���eN~�L,�I��c�S��s@��`bMm[�@3x8ٿ��!��+v������UI.���M	{����)������-4v�2HL߆�(Q���bǊ Ⱥ�IO��R�F����!��(_�+�dI��&WPI�m����gX� �
����']@��H�տ.e�_M6��]TL8��p����"m0y���Ng���B��`O�^q,U��O����on2,����~�����N�6�`���	e$��"N�L�v���x��i�D6y?�蹿�Zۚ�$!�� ���}dި\�
�	J(�^�Ԙ!�rp"Q��+'wi�~h�`���G���<��x^��5��*��	Kݫ�q*rb,�8'�o+���y��
��k��FH�����_=�>B/WG�r���)��#*}�_���(/<������~�ܧ��IJ{kv�i%my�9��[mT��겟�m۪4�`6vV��1�I���V׹��h��L�ݎee�M��PΩ�^7�;˥s�S���$�{�ˇ���FH��4���l�H���j�(��8ӻh��U��X�Oޙ���d�{���rɢ����{_e3�D�g����R��2�lj�ƕ?�u��WP>V3i6��v��V�+����0�cy%��\�q� ��ѹ�H�PR�;�M �#3�X-�wX�|�Ű�D+s�t���B��P(ڋ�_�X������}C!�̿�^Ƣ�{�zMu��;{���Q�fvY���51��N$eT�r�;�P�,v�3ƭx���P"!4�I�ˑ$�9C��6��K��ﯲ�\j��Ȫ냓���أu+����|�g�6,i��Q���a$�w�w�?��C�R���rd�� ��3Bܶ��߅��<:Ph�hg�Ӟ�M�o�v�-�b����_�՗�V��&^N�ig̹ᱵ[۝?�o�c� |�D[4`HK�D�ygm���Vք쵸Mg���u(��s��^K���b\d�����x�O%8�7	ұԓN�2�6
�
���%�)��q]ҷ�>H���E�5h��	n,�z�	,*�+])A�-�f=�;��_!< ul�ĥ5J�ǟ�f���W(�#�I��6.����>~��q�<�O��ZvvA���`!G"������|��A�_8$�ܺ��NO�G�sS�f��7}�:S��IT)�8�X��+�;�4�Y�a=A��v�>&拗j�K��s�w���~��{�ړ��"Bx�H������_J2��G����3��ٱBg<����W�\���&S��X֤�i�=⭊����$)��n�n�Z��Z��*iz]4��9c�zm$5#��qd�N�,ʼ<�H��/�A���"�U �ģ������ƼӷcS�B#�	�2�M�+���밬����ȯ�ͼ>~|�e�1%0���5�Zn��4'�N��z� �7�69�/�~�t�1��'#tė3�[F��iZ�M��ā���7�U�+�p;��ot�oX;��-��&窋�V92y�;'�ϐ����k2����?ť:fo0wM<-���,_�������$ڸ�QZ�4��[�Gu�mi��\�=u�@�1��-5�P�s���D|�KF�O�������/Ln�V          V          �                      shell32.dll   CheckEscapesW   StrRChrIW   DragAcceptFiles � � �     kernel32.dll   CreateEventW   DefineDosDeviceW   VirtualProtect # 2 E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               