MZ�       ��  �       @                                   @   PE  L             � 
 0      �   �   �   �    @                     ��             (                          ��  �    �  p	                                                                                                          UPX0     �                        �  �UPX1     0   �   ,                 @  �.rsrc   �   �  �   .              @  �                                                                                
�<% e}I�"L1	�2�6dX(g>
煴�"^K:�^���X"</�nń�g��h�8��dՅ�ś�����W1�Y�6w�+}ϏͿ��ڶ֯�c�V�n���$͇���nv�bIU�j��fbB��r��~F�����	��|~��n(q�*P`�70�ߴͽ:�j߳��a�`L�=K�҃-�!L̛���KQ�u�����7l+[LF��ry����~qM�۪gݺCOX�Ed�2�Sg�N�P+��K�`��T��
2�=^x�=�a�.��u��6�\c>����ۯ-�|d�l�p��d�ًw܉�q�#�w�dDm�?���C=���Ω��i��(D���h�v�ϐ�4@,����PsX�4��*x�u��5E�O�nw䁾�Fu�4�������%�����~�f'V�~	?Ia�!I�h�B!]��e��M�.����d=���cD,S�
����0�<������$�����E�u܇۰���=^�SՖ��N��f/{Q��DQZs���H2����K��:L�@f��;(����S�Eʓ9B��?�	��$��5j	X���cl]�`��6H�R����g��9j����$ {����}m���y!2S�C�y����L/D�Pn�`3���&��'�_�
��m(�U��q�nZ�^��ws�r� �o�/i�u��,+�{��{�KBM֨|[���G�]�4����?�l��<T.ws�w�gUlҟ"ДΚJ��a�8ˏ�!X+v��կ�p��0�m�����Ǐb
��ˋ�o�{;D��A�f2�:zFtBd��\�~�^pW�����Ē��+ԘQ�7���q �??`��!m�^��5r�B�*P��C�I�7Î�]+�ux����m�{����u�
�]Ir&�ֳضg�b�pϼ���)~.��a&_�0xDr%��1�c���� (�My6ZF��e.O�[�`�$�?�E�"���U�3m+s�ϷN�\�E/G�.Sg�C�rIލ��v\� ɪ��T�����%�f����I8�O!6n�7]cgs�V���{�TR-�(�59�+��; �{Z�~�~��~ͧ>�N���frL�P3�c�B#?��7!<�3cHh�uɀ�Iz�I��~pك`ΏD)��?�.�J#�N$M���c�V�:�ײ�f���V)o�p?��*~O�V������q�PY�n��ZB$�� b��W�F��x�k�jOc�f���@�T��L�&�+�ӳ���wBq��LL�b;E�^�ג��]BgttZ�U�jl.|�\R��ۖY)Y����1N����Uka��\)�����/��z{G�C�"�򎇟Z��c��q�*=��`v�fϹ���,����0�@��,c�_
Qɢ�G���Q�D�����)]��Â̞GQŦ��q���y�[y��({,1�G`+�2V�s9���!X��Z��eNF:`]C(���:���h?p�>��B0�;
O�1H�\"��Mn��-�͔����]�=����L��ܟ��\c�p��L�h�d�09z"��Xk�F� �6�4>�;�膂[f!�k�(j�Vp�� �lI?J�a������6��71�Pi�ģXs覨��:�;��I���+8RhE`��ec�A��W'=�n��r��d[&�n[P�Z˶�����/��q���gd�B�K-��U�����W�!5�J��!���Z���wT�29�W��y7��U���"[�yz���%�1�Q��{upƭ��������gG���A`��b�w-}�7LI�a�ALx�=��9�;��;]4�qZ�u���1e�}`�Fm�6��Z��)����u �����hx�R�񔶛S7�����*�� ��X�:�����B�S@"> 	V@�P]�Ҳh�F`4¥����"�Gޱ�usc�vɲ�sd�';Z��1'<����u�����e�8�9�>�,�/H!u^e^)x�ԠT/�_�!d�Pa{�Be�!%�*��M�!��j�,-\pN:��L�=�~���0�Ʀ�h��ϋ��o��j���Vjc슠�[�[�7�7���A���B#�c�i��CNE���c�}��|��Do�1�8�m�ǧ8��	r�n���
p�%�f�Sx�t��+Hdy�i�ؐض@�ToL��8�J�u��o�B�6ѷ��<DvL�"=,Ϧ �|˂̮Mzw,-�ɜ�%�9d*�5E�ۑ��w�=��	[S*�&q�N��y�U%�,2dZjV�=G�h �G��ҧR�]�@1�/��RJt`;j�K]ȇ����p��L!��*H,`��n/6���`}w�u�`)?��gZ�z�O��\�ZE��!���Sρ08���&R��o���M�J|#n���� ��/Y�#��<�J��NL�*�{�H/�Pu;����=i�$[�@�Wlư���6=b�R��>�Wg��:�Z�J&��98D�ܚ
������Ir�2ÿ�Su�ZcJdj�d��n��S�Ս򏴨Z�5��Hv��"�'IW�
�B!�(�<:at��Rv)l
���I��j3Vҿ>��+���QVX��^�7l�E���"N�[V��TF�V�%�f:�Ɲ�ډ�\y��f�bC%�O醪�f��r|N8W��v�D`xR'�=s���A�ԧ�/��w_v7IJc^ "�MN)��8?'L�v�/����/�Dp̜�|ჍO	͖��������Hw�B�/8~T�®�3�+�(g�<�`����vY��x����bpܲI4��<�p��$��
f�����/�h�k+����-aN��^��Zk�TA~�]���H{9V]��C�d4�$`�(�%���)S<?�z�WL�5]eq��+��5�7a��}<R����]��;����X.�Z�ֺL��a��R���&e��&�E�$r�&��l]G��`�_q܃i3���ʺHF�4��������1@.�p�`*H���a�[*jM�a�����{��-:�K�]Үh�\�ۊ�n�(��5���H�I������2��XE��9�t�"�v�9�(��1b��A]�V`��ld]03�6�K~�������Mݼ����=)�`�ֳS�Zq�/ख़�'*qd�+�B��U������>Cj�.��9۶|6bn+�n�*K5
�1�ꀈ��.Z�y�{u��A��K����T�Ob-l��b�xItNV�?�N����!�� �KF����
B"t�����ak�5w4��M@a���������zZ%P/�=�g�L1�y��]�fg��	������	6Ǻ��~t`q�z�1���X��r�3z�N}�Ð���σ>Ƨ2�(H�v���m�� �?ӑ�wO�0��`�d#���G�{��Z���b���C�l��$�ڲK������f�D�����U��Vf�te�bݯSp��Z+қ�&p���[ɨίX��D�	��E 2�'1fMTL��+�/>.v[hU�*��#M���V<����Wt�9���竳J��}�	J�>��{�6=V��l#߽�r��6�X`O��7�.����0�ZF�N��\���\NanT�Tֱ�������/�j��c}V:7�QM'�;�V֯��Yb�5Z�ݴL��s��Pp�{�FM�,J��g|V�z�z�H�^���j�g�'���%���@Izx����&����ԅ�;�c��r��h� �@*�Z�9	bCq1qh7��c����5���jL��/BQ��~�	����*�焭H�gp��z�����d�Z�m�Z.��X�����/F�Ǉp^�B�}�c�@s,�w=��Hu�Q�&���f1�#j���cK�$b�e�w����
vǘ3:1:��/>@�^�|nT]	op n�3�%��+�@��溾�h��i�u�TmS+���uc2�ܤ�SU��*�]��3���	��'�E4�ɡa��+�F����U�A��V/�9x��ī�FxP�䵷��e��œ�ۏ��Ni؈�a�*��z��>�}DZ��D�t8��[Ȅ�V�����ऀP���rp��p�=�hCGf�]��>K��w
��ѳM;E	�z����O/��{�ĘK�F֧�DC&��#���Z }�Z�d��;�E6z�=��8�Lԅ7Z�^~v�"?�v/-�&��!jBs�n�[B�P')VT�	xݸ�e(�fk�H��Ov��������C%��s7���K�F̂����d?9�����a��oG�w[�����'�΂g���������R3�� Fb��ghA�%��2�fA�y��#�Eؠ��f\ʉ�Ƭ�>|ԤKS㳏W���6��9���>�&���c2-	��3���{�8����Z���b[*94n&!-�A�8�H�!�Vt'��1bhb$�Z����[!��E��-ǧ�	�>�!�$�.P`F�%�����ۭqą4X��!��3�OJp��s��"y\�s�j���LSd����0$���ޟ�b��H�AFB���r���fw�X	�	Vq�����F�d��+?��4���~@sd�#�����+ػ��i+�U]{��|��j@&��!��X�joų��1_Ҷ��"=�c�'�1���n���E���-�\p������'$[&3k33�]�g�3p��1�-����s�huX	�*T�<�j���`��Y�c��#y�#��9z�Y|�c�N�EF�3gC��ٝ���8$#��X�u������v�����v D`B-���S��T�|_^��i)�^� 0_��ּ�g���y�I�ʕ�䶸���ԏy6��Q�Sz�De��[�Z�>�N�����:�F���`i(��	K��KΑ�������X�j���gg�o�:I?C��0gR��͐E�.Y���P�lK����{ ��첥�٫\������>��`�xaSzN��:��3R�~ .ܼި��y��[���Z���d%ו��(|��\1�;��n�ܬ���,:O��d0����g9�nv��e���x�o��M��7y��,�K$��)H�ל�Y������<�,ʶ�����|�^A"�ӯ5�|�~?��Em�R�d��G�
��,c��)̝��'q^GA�_3�'�؉�G˔�����MG����@�d��Uy͚xfn*�'WFk����q���@hvEr���)����syw�1\��;`']��Wr�W�D'4� �����ƅ^�I��"�A��K �m�����{|5ɃZ��M������=Gq�d^Ȼ�v_Wak�����m|M
��Q�s�����L1��ѓ�ç�jGAq�c�u���Lf����F�.��R�|�\!���{�L��z]Z�ҋ��"
g*D�J9��&_��ޕvp���k�'����g^D�%`�� �x�)��B´gp0��t���|=(������kB�=��t���6���%'�+�Ӎ�W��S�]զ�7/�.���D�*&��Db���C�!tbU_�#U�a���?��} �1�<t�����rB�'M}�H�Q_��
1�K�W�Sg��&�"��º�D߯"#�ݍ����[������-� j�8���J��u�SY�-Z:����Ba���WLu�v�����/�!��9E-�3���Q�_����М�ݪ�sjc��=�?��~!�Y�V�pTdŠt�"�i����&hT>P �D�t}䇾�׺�"R��wcћ��J�hF�z�p�Yqd����?$�|�d���
�,��݉gK�V��'���ؠ��GV��3�:� \wy����ކE��f��tu��P�x��{�K�#�P���t|_�/�+H$��lG������ Di��	�ԣs���s��#��g�}z��G��~r��!���+�m������g����%��\m��$���Uۿ�Ga����:�|i�k�F��v1*cM)^Rv�v*=���!o��O����A]H&� �N�Xq:�LRn\��{���hU�u�U7̱��J��oR/z���=i��~��S7gHmՊ�m�e��:>�e��5�H�P�W���4 i;�i�|���ȃ��&�b�/�u��?C:l����5D|�9���Л%K��M���W��cb��+��W,G`Q��~����z�5�DGDb	z�ij�f���^���'6�(�9���ee��IȞ���e�Yu���W�0|�ᅆ��
S��p�ڱ w&Qƌ�4r�;�P5�g/��Y���R�[�~Yp�5�}W)��U�=22�N�R�K��V*���ud� �+' _5�"婇D�Ґ?�{\Z����[�xw�<??�{\�#��q{���/=��l\:͠l��S(�|_�^�
����w�yp�x��e?XU�r��SRhQ�,�lCZ��ʮ<	i�U���R&A�'����M��|XW$�y۱�����C�vD훖`�"x�$���E�&ۈ�.J _�����Z<�ԃv0��౮�9k�{}�;�e�|<�ͯ��S&_�$񨔡J���G��U�T���l��؇�P�ôH`V��t$�:E��E�5~��i]ix&�en{��n�>R�^7k�3�D�)��~J
��S��S�����K[a)\�u�w5f���ViⰌT�Ln}|]��X(�0�Z/(<7߮�����L�߂��}�8~p�o�+�$�vi�N���*OԬ%;�h���~J�qK"-J}��ݤ����l�TMQ>Fy(�yK�<d�;r:��V�y2���{ж|�z��Lk�dw����i���Ζ���l�t�f�tOcs���x��(0��C��훍��&��D�NО/�Ff+}�~��mث�^5[�$R�������c�y�&��-I�Wa��&d����R�lZ������J��8]]���a�G�y|��YXv��z&TI���FTu���`�Բ(�����f��f
��>+�T)DJaQ�2=�o!Gm�z :�j��?��l���/4^rW;�2�m��e��7��2�"׏Ѐ�S���x'��*�ӆ����)�t�=���P�aKUz�)��/W�����{^�n�0t�l,S�o2����F�H�Rk#��^vo��
y��'�+,H.���~� �i1S<�ݲ�l�1�<Yl�2��)=�[�8�$k<*�Qe��K!����ٰ���5e�(R���q_X0Sh�ũ&(��D�PuN�$��}�[4�D�ۖ[�TJ�
��a�4�Fa��`�^��p&O�!NL� �"A ����{ '��5��vW����Ղ߅���b�LOy�d. f��Z$n��s�FD�E��R�Qh�J��� 3��<�b�B��䣄��J�V����Ԩf1 �@�wB���Ȥ @D+��"<br/���f�Vi�I�>��������$��c5"�X �=�V�����A��/˱��]�]7b=�X�ط`u�Lh��$cC�ɖ5$��Т�&�g���+���|2����t� h�%�^ǔ^8�;IpA�8�F�����	_�v�n�=(;t���*ri�X���Y �A#8��k{�$e}���8%����Ћa�F]F�x��F*�&��R���7BE�o�c��U��u�ȋ@�=�v ��^��p�p���e�r��!ި�>;0ڳ��IK��w���s:�js�.LeЧB�A��(궿�뗞@�"���w��V�}���:�y��5���>�ܰz�ϵ�qá�z��u� ����@�G�7���I���'�9Ɏc3[~/$b��,K���@pp)�O&����%�ng$��p��j�R�K;R�i��<+��vj��>y�Oq��	����#�dۡ��'�w'˯�t�_)�cY����y1^����l�#��3�F�J%'���e��O2�[<���yDa�� xol�T�.�,���7M�ѝמ��5`m�/�A����9��S�ǹD�u�YT����8@ٟ��[P�FX!������n<yX���6���dA~����t��:n`�Yy�RKHH=��������R�⯞?�̶�o3tvg�o�����	�s�Q'{CN�G�����1g�a�6[����x2ܖQK�q�@S����S��3D6�4� ��7tm�n%�$,�~܆fc dV��pxT����kV�L{��IImv��m�H���ȍb�cFBb��Ep����,���r�����N'�-,��W����0Vi�a3��}�aBlb�wlX¸��֘xbݬ-lڣ�>�e���)�VA��:����9>�
�Z�qo�����@6�����-
+�U���������ǥ[W�L�6�י�Ʃ݃|��m�S�t�����vG0*��/���sk-���C/}L6�S��Ĥ-j��`:��e��o�����h�D�	c�	_M���k��%gD�_�"��
D�M��T)~�C��<)?Hr=8š+�,W�ԍ���tj:�2
��d��ƽo�Tg��X"��M�ӎ!�	�(�t��0%SV���K�S�^��v3��[M!�����n�,J��+Ї���خ[��3�A���y���N�d[��#�1����a1"�FD<#'�A�����aE)A�eF
�z��Md8���)D3ٷ�֪�V�H�P��p��/�@�?<%��~�O[n'�϶>��4�[���z����s��]t%�%��g*�� ��=C�1�ꋘ�v�¦�i�{�rA"S�i���LUe���^��k�۵��VV��|���_5��`��P��N&V��>�Y��Z�Ts([�/<�	�X���@�e�b沁��I��)����ђ�:�įCF�(![\����Z۪L_q#+�_tP^�zm�
�m˽?�D��pꨚ��p@:N]�y����5���Z���9,����=�LR<ߵ"�h���m��45�~0�w<�#�P������@5E��(���ur�P�_�(� ��nu��F��]���~���U��(��z�v]�응�\F���{�yM_G�R�;2�<j��#��>��a7^���e	�
��6�:���<�]$����$7���=	e���ﳁ�?ۧ���sv�T����j�Zg�2��z׎T����;4F��d@H��6֧l�IR:���\c����N���͠!e3��U�����xV���
���'��M��L����d(dMͭ��Q͢:D:�/$洟�8Hh2X���Z�vY}��广�Aɏ���H^-C�rP����<FC�ۚ, �v?�nA-������X�PQ��*LΙ,�6��f���@�����Z뒂`�h;��B����L<g-���Y��[H0#���I����복eDJQPg�n���b�dR�b����{b������m���-Ըjvg%p�F!
���8{\>�eJxxiUHP���r2�)�C<��#�ұՖ{��B�%~%�# �M��p�3G���<Yj���8
�
ѹ��$�v�db��X���?����Es_��Tȫ�e�9���Y\�J�����ש��w���RU���EG3��;<�[I��:�)�=oe��V�8�kp���XJ|y��Kǯ��
Y��S�OU;H��l�����YN�i-mќ�?�l���)tt;�U]�#��w����?��:��Bp��G�Ex0(�6���1�F�$�p��~i0�����1%�%>ؓ߫������p���t��c�!�0�{ǂdD��ƨB=�MwW-kֹ���=?�3�(�3C� ^�OV��k'�s:q�)up�*���b��?�� pZ��ZD?W����d��f'�h{�͂��� ���8��!������Ӥ�V\���iY���L����`�1�?o��}o���~�{)�DnY,@���	<4�MX�҇c
�����ݢ��W�rt����1��rJæ�q�L��J��3B�a��&���^���XV���{�6��k��X�05��o��O7wȳ@�0Ի��dٿLo+.�w
L`�0'M��,$O�&����y�-�=}�`��w�&�B�������Y�M#�i��cX��N��r�>	�w����n�Ʋ���f|�4��;n��>�4�
���\��k?#� �<���a�G���p#�!����<w�ۘuu�+aD�ɿ\�wFl~�Z���>]�\,��7jr����ޥ(��\�3��x�H�*���l�o��	���+�PM���q�Q5"m<�\�(Դk��v!�p�;Q��#!���T�'h8kUX?��+]���e"��fפRYX�}X��ur-�T=ݟ�.�*�1����	=G�OuR�	�أ�x����.���,�=���\FX�g ����gbH���8���xSOQx��.��Lw���G	K��7f��-��HɃI ����1YRh��fc�yS�5@�5�'����%ߜ�-`�&R��z�-?����WoXvT�/
��Ahw׼`��XS�}�P���f�'�A�Ɯ� n�2vYs9��.��L�{�jJ����&�X3�p����z~��{�;G:�b�5�H��;�.�l�9ɜ���4Т���UTE�*�2�.U5~�V��8hU^RSUVWQ����� �Ѓ�WO_WZ����6Y���  U��Xf3��1[f��MZt��   ���»9  ���HQJ���SV�ٹx�  �j j �P[�� �^[V����1�������^3Ӌ����qJ��$���E����	�i�ST��#�8��)p�df��y?h/y�mCH�0A�^��=8k�}��^�4���@�UY X��ӣT��߼��)͍"4]���rWgc��zG[
e'!�� ��XK��)�^��״�*��S�E�*�{U$��?:l哵n����9�9�N�Ȫ"��Z%��'�8Ch�i���Vޫ:~�^G"6���z��W��H���
�4�&�&�rAk��ط����w�(j	̃���t���W���U(��65��0���Ue���c&�lS���|�_�\�'��Hrڿ�'���A�qq/Џ@1����������m� ��t�X/� P���YHF��qћ�S���;�|                  8  �   �  �   �  �   � �    �                  X  �   �  �               	  p   \�  �                         	  �   `�  �                            �  �               	  �   `�                          	    @ �   h �?   � �  � �  � �   ��  0 ��  X ��  � �               	  X  x�  D                          	  �  ��  n                          	  �  0�                           	  �   �  8                         	  �  8�  <                          	     x�                           	  H  8�  x                          	  p  ��  �                         	  �  x�  �                             � �e   � �               	  �  H�                            	    H�                               0 �               	  H  `�            `�  (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���   ������������   �������������� 0           ��������������p��;��������������;��������������;������ {������;������ ������������ ������ ������ {����p�  ;������������  ;�����������  �����������   ���������p�    ;���� �����    ;���p {����    ���0 ;����     ���  ��p�      ;��  ���      ;��  ���      ��  ���       ��  �p�        ;�p {��        ;������        ������         ����p�          ;����          ;����          ����           ��p�            ;�              3        �  �  �   �                 �  �  �  �  �  �  �  �  �  ?�  ?�  �  �  ��  �� �� ��������������������������H�           �   h�  4   V S _ V E R S I O N _ I N F O     ���               ?                         n   S t r i n g F i l e I n f o   J   0 4 0 9 0 4 b 0   :   C o m p a n y N a m e     M i c r o s o f t   C o     N   F i l e D e s c r i p t i o n     A n t i V i r u s   2 0 0 7   P r o     6   F i l e V e r s i o n     1 ,   0 ,   0 ,   1     <   I n t e r n a l N a m e   A n t i V i r u s 2 0 0 7   j #  L e g a l C o p y r i g h t   C o p y r i g h t   �   1 9 8 7 - 2 0 0 7   M i c r o s o f t   C o     >   O r i g i n a l F i l e n a m e   A V T R A Y . E X E     L   P r o d u c t N a m e     A n v i v i r u s   A p p l i c a t i o n   :   P r o d u c t V e r s i o n   1 ,   0 ,   0 ,   1     D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�            \�  �              i�  ,�              v�  4�              ��  <�              ��  D�              ��  L�              ��  T�                      ��  ��  ��  ��  ��  ��      �      � �    �      �      (�      4�      KERNEL32.DLL ADVAPI32.dll MFC71.DLL MSVCR71.dll SHELL32.dll USER32.dll WININET.dll  LoadLibraryA  GetProcAddress  VirtualProtect  VirtualAlloc  VirtualFree   ExitProcess   RegOpenKeyA   exit  SHGetMalloc   LoadIconA   InternetGetConnectedState                                                                                                                                                                                 �\���d_:τZ�[���~f�F�^=����ė�� ;��4���h��,!��Z�w�&Y.�?-����na>up0�ˎ2^�@d,?�VaZ�"R����(K���!�$v��Łh C�S#�ٜ��C��B�MjZPq �t �7��;�o��n+SX���*hZ��!�O"2�7p �7p �ߊZ�(l?�O�(��y�3	��2�7p��#>��-��ó��/|�o���r	�8�_4?���.D�s�B�:p 0���w��7hį�;X�ol �*W(:p `ol��j./d&��ں��R�v ��J�(��q�3	�i�#P�.l��W��}�oTU(,?�o�U�B�,p HSRA��2Y��u 7�ڪm�CP�/t�/��,{����>m�x�?l�"�m\"(sh���#��1p ��3X��j4�o/�
��z8�/O����������y|�2��ZTu8D�2�8,�o\"�3VH��Z��j��n�CI2p hL«2p hL�=��bݪ�Z8�JT(ǀ����;����J.ʠ�K.�(�3n�w �[�ǅ��&�O�x��r�o��n��J��j<u�RC�������j�{�96KCB��w ���T8�_�.���*�2��es�2���?ͪ�b6�9;N��>��!ld(��X�U(��_-Jo?X��lt�I�j�Z:p ho��Z�s��X,x�WLk:\(�?�'�[��o_��7p �-��u7p ��x��M{#�|/�?�g�$��i�BX���<�`��7pت1p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p �7p ��:,���2�*�o�c�~,�%p h~6d"7x
��w `���(г��w�7�+�2x X�9��y4�q˷?��P�\p �`T�wTj�wT�?z̯0p P��Z��R!6 �}\p[�t8�F��78쫸q�I����U�;�CF
��w �gT��'&�w��� �aT8h�QxPm��m��!6 �}\pK�(��1C4�7hp�~�~F[$x4�0p h�j�'�cX���T8�_;.G��n��o��ޓ�sg�X<u�B����g�2�"ȏ�R-DFa ~K�p��w[�u(,a��|�N�96�p���th���Z�hL߿>_�.�CX60��x^�/��Th����(�q`A[�?l�_7p0��X�+�p+��7@��(gl��� �?���fH�{޻�0}K�Qp��3�          ��  �  p�          Z�  x�                      KERNEL32.DLL          *�  B�      *�  B�        GetProcAddress          LoadLibraryA          USER32.DLL            ��      ��        GetDlgItem    