%PDF-1.6%����
17 0 obj<</Linearized 1/L 9915/O 23/E 5149/N 1/T 9528/H [ 716 170]>>endobj                     
xref
17 21
0000000016 00000 n
0000001053 00000 n
0000001202 00000 n
0000001241 00000 n
0000001282 00000 n
0000001326 00000 n
0000004085 00000 n
0000004305 00000 n
0000004367 00000 n
0000004397 00000 n
0000004430 00000 n
0000004466 00000 n
0000004522 00000 n
0000004556 00000 n
0000004691 00000 n
0000005002 00000 n
0000005036 00000 n
0000005092 00000 n
0000005113 00000 n
0000000886 00000 n
0000000716 00000 n
trailer
<</Size 38/Prev 9517/XRefStm 886/Root 18 0 R/Info 12 0 R/ID[<0583B53D49A95642808482B87A2E0F38><8DE2875640EBB8459E7C623740BAA060>]>>
startxref
0
%%EOF
  
37 0 obj<</Length 85/C 89/Filter/FlateDecode/I 111/S 36>>stream
x�b``d``�` �lL������bQFƪM<�x>(3\(R�e2``� Q��� \��Í�a`P�]` �
B
endstreamendobj36 0 obj<</Length 20/Filter/FlateDecode/W[1 1 1]/Index[13 4]/DecodeParms<</Columns 3/Predictor 12>>/Size 17/Type/XRef>>stream
x�bbbd`b``�a�   � 
endstreamendobj18 0 obj<</MarkInfo<</Marked true>>/Names 19 0 R/Metadata 3 0 R/PieceInfo 4 0 R/Pages 2 0 R/StructTreeRoot 13 0 R/Type/Catalog/Lang(en-us)>>endobj19 0 obj<</JavaScript 20 0 R>>endobj20 0 obj<</Names[(main)21 0 R]>>endobj21 0 obj<</S/JavaScript/JS 22 0 R>>endobj22 0 obj<</Length 2686/Filter[/FlateDecode]>>stream
H��Wۮ����A_]m̓g�Ǡ8oEQ�h�HY�)��E;���h+�H.޾������~��������}�~��h��$kl���`��$g"|z�w��������������������+^�7�'����Йp1���L�&�	Ʉބ��ߍ6?��H>G��&�L�R�2�3)Cxɛ�O�$�9�4�w10;�q��h\2�7n0�j��⮦�L7�;<
��Γ)`�f0߅3~�c�-x�76�A]�����Bl׼�1��=k��������Ŧ+)�ca��X�y=녀}A5CMS�5ʌ$���֍���A�M85���K�y{r���J���j¿h.ǉ�ɺvܲ����{�a=@�
�-�Aw�3�;R6\�/ȡ\G���d�L;�8���K<f�^�.�	�W�U Q�1,���&`ԕw� W��������cf�#����� 	?k�.�0a�v} M=Sۄ
��K.�ڱ�K��&��2�K���hp2<\����<
�S�u9[J�B�W
�u�����3�~�dC����o��/Xkf�Ϫ훂���-Yb��� x���!��ؔ��g�G_��E�U�r|+P���4Bn��b�t%�/�����9�J	
?��`&ێ��Rڒ���#�=_q�WJ!�r~���X>�qn��Hų���u�AZܶ�^�q�_�߆��������^���{xK��W�1Y����5-�5p�uudъYR�+b�p������1�`�Wl��N�O��	�xH���ؐC�k���܋]z�m?�h��:����Q�-g�[n�o�VB����><���0,@S �{��3��;���б��sW��8CF�0_ *�	p���i�y�σ��|討POFCPو�aNA�f��><�|=	O���Q�?������T�.����D��˰Vv�^����6�}9N�w�u�m��J�o�i�h�wS&F���gE
���Z~�d��{��p�L3�V�Eͺ\
m`�Dlj��������S�qȍ���6�{��z�L��Oeg��8�7�n�rFF*x��c��;�\��������|>1r�$�}�0p�-Ϟ�rv�S�����J�Uw�JNûa���˟*l.�[�p"6����,ɱ:](o׻S��ݷZ֢��X��J������[k�O�� ���rh���>��o�c��Li�#抆X�؁r��p�R��>ۼ�)���(Ǒ�^~~!���n����>x����K�*��ą_G�5��-�y�^h�����A�^v$���>��-r�xi�a�aW�6;K2����q���ʺ��zi���Z���� �wm����l?p��r��ګS�ru瀿*�hgI/*�����0h�lyl����@=��50���μ������?ug����y�j%^����?��q6�-�}Qc���XC���.��9P���.�D�G�yx#�)估�vέd^V�ڸ`kP�ȫ�8��d�|!�P��Z�ף������~�E���6�)~)o(���w���%����s�Ѽ��+�����𕿴�9��Ty8	z5�AQ/�}ޕ7X���p��g�s����T��Ϸ�GʥG������`�{��R_����Gk疜��_��YYO���ڭq.�R�yi�93�h��?��N�_�̫�S����o���E�g��zڟ���z!a;�wa�;�����Z�j}�^�_��MP�b?���޲��R��r$��E[�)�?O�׆?�zᄵ�ϒ�����K���lr�>g�ޖڪ��m������8����Q����}���s�������!�ug��?�멐��������ϟ����~L�i*<R.��㹼���$�5�E���dg)�N��l�Z�]#.������x�:%գ�9Q/�8m�#Ʀ��j1�>0_�3-<��p6���l���9W򻺟�r��>����Rk~�x<�>����y��O�)��0�h�1)f�zI<T�]�U����#���v~i�!W�������Kʫl?���|��wmސ򏶏�x���d�рg�?<�1f����K�ש�iW��i�i��)>��?o�#�_;WJ6�:;����/����\s7~�Y۽��*��9�_��:;����]��}j�� ���5
�s��{J�[�\�\��S�#�˧�����+������i���&�V�O�mYl��g<�хrf�CG�F�O����1r����u��	�7���O��q�9��(�N��8i"aB��MG��V����3�����>�~�t�c���_�����c�ث�n{{����?��n?�c��N�[����Ɲ�-��]1�"G��]����t�r��S��<�8�>�&g�3O5���� �m���^=q�6<�dzA&�}�Y@��&�9ƶ�r��z���Q�ۇc\=ѻ��&N��fdl��=�'1��~�����������V����� ��#k�y�����ë�Fk}����l��J�����ˢo5��=���{�4#T��덏h�\4�7|�pr&R���>��4ȩ����s�ce+�����	�s5	���PW��hg�P��\��3����,�q4������C0��K��]>�����<�k����~���� �
endstreamendobj23 0 obj<</CropBox[0.0 0.0 612.0 792.0]/Parent 2 0 R/Contents 24 0 R/Rotate 0/PieceInfo 32 0 R/MediaBox[0.0 0.0 612.0 792.0]/Resources<</XObject<</Fm0 31 0 R>>>>/Type/Page/LastModified(D:20081110184212+01'00')>>endobj24 0 obj<</Length 12>>stream
q
/Fm0 Do
Q

endstreamendobj25 0 obj(DefaultFlow)endobj26 0 obj<</Flow 25 0 R>>endobj27 0 obj(D:20081110174212Z)endobj28 0 obj<</Private 26 0 R/LastModified 27 0 R>>endobj29 0 obj<</PDFWP 28 0 R>>endobj30 0 obj<</Subtype/Image/Length 1/Name/X/ImageMask true/BitsPerComponent 1/Width 1/Height 1/Type/XObject>>stream
�
endstreamendobj31 0 obj<</Subtype/Form/Length 49/Filter/FlateDecode/PieceInfo 29 0 R/Matrix[1.0 0.0 0.0 1.0 0.0 0.0]/Resources<</XObject<</Im0 30 0 R>>/ProcSet[/PDF/ImageB]>>/Type/XObject/BBox[108.0 72.0 504.0 720.0]/LastModified 27 0 R/FormType 1>>stream
H�*�2T0 BCCs#��\.}�\�|�@�B����	P� U � z�}
endstreamendobj32 0 obj<</PDFWP 33 0 R>>endobj33 0 obj<</Private 34 0 R/LastModified 35 0 R>>endobj34 0 obj<<>>endobj35 0 obj(D:20081110174212Z)endobj1 0 obj<</First 23/Length 105/Filter/FlateDecode/N 4/Type/ObjStm>>stream
x�24V0P04Q06V04U03S04S�4U����	(�T����&��������A��(���.�ɥ��ypf0&P�E� ��`}G�@� ��"8
endstreamendobj2 0 obj<</Count 1/Type/Pages/Kids[23 0 R]>>endobj3 0 obj<</Subtype/XML/Length 3493/Type/Metadata>>stream
<?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 4.0-c316 44.253921, Sun Oct 01 2006 17:14:39">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:xap="http://ns.adobe.com/xap/1.0/">
         <xap:ModifyDate>2008-11-10T18:52:28+01:00</xap:ModifyDate>
         <xap:CreateDate>2008-11-10T18:42:11+01:00</xap:CreateDate>
         <xap:MetadataDate>2008-11-10T18:52:28+01:00</xap:MetadataDate>
         <xap:CreatorTool>Acrobat Editor 8.0</xap:CreatorTool>
      </rdf:Description>
      <rdf:Description rdf:about=""
            xmlns:dc="http://purl.org/dc/elements/1.1/">
         <dc:format>application/pdf</dc:format>
         <dc:title>
            <rdf:Alt>
               <rdf:li xml:lang="x-default">Untitled</rdf:li>
            </rdf:Alt>
         </dc:title>
      </rdf:Description>
      <rdf:Description rdf:about=""
            xmlns:xapMM="http://ns.adobe.com/xap/1.0/mm/">
         <xapMM:DocumentID>uuid:efd452b0-84f5-4a3e-9779-5c07996877cf</xapMM:DocumentID>
         <xapMM:InstanceID>uuid:fd0f56a7-209b-4f91-9a7e-208b9fadee64</xapMM:InstanceID>
      </rdf:Description>
      <rdf:Description rdf:about=""
            xmlns:pdf="http://ns.adobe.com/pdf/1.3/">
         <pdf:Producer>Adobe Acrobat 8.1.0</pdf:Producer>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>
endstreamendobj4 0 obj<</PDFWP 5 0 R>>endobj5 0 obj<</Private 6 0 R/LastModified 7 0 R>>endobj6 0 obj<</Version[1 0]/Flows 8 0 R/MasterPages 9 0 R>>endobj7 0 obj(D:20081110174212Z)endobj8 0 obj<</Names[25 0 R 10 0 R]>>endobj9 0 obj<<>>endobj10 0 obj<</F 11 0 R/Name 25 0 R/Type/Flow>>endobj11 0 obj<</F 10 0 R/N 11 0 R/O 31 0 R/P 23 0 R/V 11 0 R/Type/ContentRegion>>endobj12 0 obj<</CreationDate(D:20081110184211+01'00')/Creator(Acrobat Editor 8.0)/Producer(Adobe Acrobat 8.1.0)/ModDate(D:20081110185228+01'00')/Title(Untitled)>>endobjxref
0 17
0000000000 65535 f
0000005149 00000 n
0000005348 00000 n
0000005400 00000 n
0000008970 00000 n
0000009002 00000 n
0000009055 00000 n
0000009118 00000 n
0000009153 00000 n
0000009194 00000 n
0000009214 00000 n
0000009266 00000 n
0000009351 00000 n
0000000000 65535 f
0000000000 65535 f
0000000000 65535 f
0000000000 65535 f
trailer
<</Size 17>>
startxref
116
%%EOF
